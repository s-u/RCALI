%!PS-Adobe-2.0 EPSF-2.0
%%Title: integral_geom_4.eps
%%Creator: fig2dev Version 3.2 Patchlevel 3c
%%CreationDate: Mon Sep 29 10:04:11 2003
%%For: kieu@tulipier ()
%%BoundingBox: 0 0 495 350
%%Magnification: 1.0000
%%EndComments
/$F2psDict 200 dict def
$F2psDict begin
$F2psDict /mtrx matrix put
/col-1 {0 setgray} bind def
/col0 {0.000 0.000 0.000 srgb} bind def
/col1 {0.000 0.000 1.000 srgb} bind def
/col2 {0.000 1.000 0.000 srgb} bind def
/col3 {0.000 1.000 1.000 srgb} bind def
/col4 {1.000 0.000 0.000 srgb} bind def
/col5 {1.000 0.000 1.000 srgb} bind def
/col6 {1.000 1.000 0.000 srgb} bind def
/col7 {1.000 1.000 1.000 srgb} bind def
/col8 {0.000 0.000 0.560 srgb} bind def
/col9 {0.000 0.000 0.690 srgb} bind def
/col10 {0.000 0.000 0.820 srgb} bind def
/col11 {0.530 0.810 1.000 srgb} bind def
/col12 {0.000 0.560 0.000 srgb} bind def
/col13 {0.000 0.690 0.000 srgb} bind def
/col14 {0.000 0.820 0.000 srgb} bind def
/col15 {0.000 0.560 0.560 srgb} bind def
/col16 {0.000 0.690 0.690 srgb} bind def
/col17 {0.000 0.820 0.820 srgb} bind def
/col18 {0.560 0.000 0.000 srgb} bind def
/col19 {0.690 0.000 0.000 srgb} bind def
/col20 {0.820 0.000 0.000 srgb} bind def
/col21 {0.560 0.000 0.560 srgb} bind def
/col22 {0.690 0.000 0.690 srgb} bind def
/col23 {0.820 0.000 0.820 srgb} bind def
/col24 {0.500 0.190 0.000 srgb} bind def
/col25 {0.630 0.250 0.000 srgb} bind def
/col26 {0.750 0.380 0.000 srgb} bind def
/col27 {1.000 0.500 0.500 srgb} bind def
/col28 {1.000 0.630 0.630 srgb} bind def
/col29 {1.000 0.750 0.750 srgb} bind def
/col30 {1.000 0.880 0.880 srgb} bind def
/col31 {1.000 0.840 0.000 srgb} bind def

end
save
newpath 0 350 moveto 0 0 lineto 495 0 lineto 495 350 lineto closepath clip newpath
229.0 123.0 translate
1 -1 scale

/cp {closepath} bind def
/ef {eofill} bind def
/gr {grestore} bind def
/gs {gsave} bind def
/sa {save} bind def
/rs {restore} bind def
/l {lineto} bind def
/m {moveto} bind def
/rm {rmoveto} bind def
/n {newpath} bind def
/s {stroke} bind def
/sh {show} bind def
/slc {setlinecap} bind def
/slj {setlinejoin} bind def
/slw {setlinewidth} bind def
/srgb {setrgbcolor} bind def
/rot {rotate} bind def
/sc {scale} bind def
/sd {setdash} bind def
/ff {findfont} bind def
/sf {setfont} bind def
/scf {scalefont} bind def
/sw {stringwidth} bind def
/tr {translate} bind def
/tnt {dup dup currentrgbcolor
  4 -2 roll dup 1 exch sub 3 -1 roll mul add
  4 -2 roll dup 1 exch sub 3 -1 roll mul add
  4 -2 roll dup 1 exch sub 3 -1 roll mul add srgb}
  bind def
/shd {dup dup currentrgbcolor 4 -2 roll mul 4 -2 roll mul
  4 -2 roll mul srgb} bind def
/$F2psBegin {$F2psDict begin /$F2psEnteredState save def} def
/$F2psEnd {$F2psEnteredState restore end} def

$F2psBegin
%%Page: 1 1
10 setmiterlimit
 0.06299 0.06299 sc
%
% Fig objects follow
%
% Polyline
7.500 slw
n 203 -1648 m -210 1233 l 1868 1907 l 3930 1788 l 4208 107 l 3228 -827 l
 2543 -2638 l 1553 -3583 l
 cp gs col13 1.00 shd ef gr gs col0 s gr 
% Polyline
n -540 -945 m -945 1935 l 1125 1800 l 90 990 l
 cp gs col0 s gr 
% Polyline
n -3338 -900 m -3608 765 l -2618 1710 l -1268 -225 l
 cp gs col0 s gr 
% Polyline
n 2268 -962 m 2538 -2627 l 1548 -3572 l 198 -1637 l
 cp gs col0 s gr 
% Polyline
 [60] 0 sd
n 192 -1645 m -213 1235 l 1857 1100 l 822 290 l
 cp gs col0 s gr  [] 0 sd
% Polyline
 [60] 0 sd
n 1547 -3576 m 1142 -696 l 3212 -831 l 2177 -1641 l
 cp gs col0 s gr  [] 0 sd
% Polyline
 [60] 0 sd
n 2542 -2634 m 2137 246 l 4207 111 l 3172 -699 l
 cp gs col0 s gr  [] 0 sd
% Polyline
 [60] 0 sd
n 2268 -967 m 1863 1913 l 3933 1778 l 2898 968 l
 cp gs col0 s gr  [] 0 sd
/Times-Roman ff 270.00 scf sf
-736 -982 m
gs 1 -1 sc (o) col0 sh gr
$F2psEnd
rs
