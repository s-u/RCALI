%!PS-Adobe-3.0 EPSF-3.0
%%DocumentNeededResources: font Helvetica
%%+ font Helvetica-Bold
%%+ font Helvetica-Oblique
%%+ font Helvetica-BoldOblique
%%+ font Symbol
%%Title: R Graphics Output
%%Creator: R Software
%%Pages: (atend)
%%BoundingBox: 156 279 439 563
%%EndComments
%%BeginProlog
/bp  { gs gs } def
% begin .ps.prolog
/gs  { gsave } def
/gr  { grestore } def
/ep  { showpage gr gr } def
/m   { moveto } def
/l   { lineto } def
/np  { newpath } def
/cp  { closepath } def
/f   { fill } def
/o   { stroke } def
/c   { newpath 0 360 arc } def
/r   { 3 index 3 index moveto 1 index 4 -1 roll
       lineto exch 1 index lineto lineto closepath } def
/p1  { stroke } def
/p2  { gsave bg setrgbcolor fill grestore newpath } def
/p3  { gsave bg setrgbcolor fill grestore stroke } def
/t   { 6 -2 roll moveto gsave rotate
       ps mul neg 0 2 1 roll rmoveto
       1 index stringwidth pop
       mul neg 0 rmoveto show grestore } def
/cl  { grestore gsave newpath 3 index 3 index moveto 1 index
       4 -1 roll lineto  exch 1 index lineto lineto
       closepath clip newpath } def
/rgb { setrgbcolor } def
/s   { scalefont setfont } def
/R   { /Font1 findfont } def
/B   { /Font2 findfont } def
/I   { /Font3 findfont } def
/BI  { /Font4 findfont } def
/S   { /Font5 findfont } def
1 setlinecap 1 setlinejoin
% end   .ps.prolog
%%IncludeResource: font Helvetica
/Helvetica findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font1 exch definefont pop
%%IncludeResource: font Helvetica-Bold
/Helvetica-Bold findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font2 exch definefont pop
%%IncludeResource: font Helvetica-Oblique
/Helvetica-Oblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font3 exch definefont pop
%%IncludeResource: font Helvetica-BoldOblique
/Helvetica-BoldOblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font4 exch definefont pop
%%IncludeResource: font Symbol
/Symbol findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  currentdict
  end
/Font5 exch definefont pop
%%EndProlog
%%Page: 1 1
bp
155.91 279.21 439.37 562.68 cl
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
210.94 325.29 m
429.41 325.29 l
o
np
210.94 325.29 m
210.94 318.09 l
o
np
254.64 325.29 m
254.64 318.09 l
o
np
298.33 325.29 m
298.33 318.09 l
o
np
342.02 325.29 m
342.02 318.09 l
o
np
385.72 325.29 m
385.72 318.09 l
o
np
429.41 325.29 m
429.41 318.09 l
o
/ps 12 def R 12 s
210.94 299.37 (540000) 0.50 0.00 0.00 t
298.33 299.37 (540400) 0.50 0.00 0.00 t
385.72 299.37 (540800) 0.50 0.00 0.00 t
np
201.99 334.03 m
201.99 552.50 l
o
np
201.99 334.03 m
194.79 334.03 l
o
np
201.99 377.72 m
194.79 377.72 l
o
np
201.99 421.42 m
194.79 421.42 l
o
np
201.99 465.11 m
194.79 465.11 l
o
np
201.99 508.81 m
194.79 508.81 l
o
np
201.99 552.50 m
194.79 552.50 l
o
184.71 334.03 (1794000) 0.50 0.00 90.00 t
184.71 421.42 (1794400) 0.50 0.00 90.00 t
184.71 508.81 (1794800) 0.50 0.00 90.00 t
np
201.99 325.29 m
437.93 325.29 l
437.93 561.24 l
201.99 561.24 l
201.99 325.29 l
o
201.99 325.29 437.93 561.24 cl
/bg { 1.0000 0.0000 0.0000 } def
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
  236.28 552.50 m
	 267.96 552.50 l
	 270.80 535.02 l
	 241.31 530.65 l
cp p3
/bg { 1.0000 0.0902 0.0000 } def
np
  293.52 552.50 m
	 312.97 552.50 l
	 309.91 519.73 l
	 292.43 519.73 l
	 292.65 528.47 l
cp p3
/bg { 1.0000 0.1804 0.0000 } def
np
  270.37 528.47 m
	 270.80 519.73 l
	 271.68 508.81 l
	 245.02 513.17 l
	 243.93 517.54 l
	 264.90 524.10 l
cp p3
/bg { 1.0000 0.2745 0.0000 } def
np
  267.96 552.50 m
	 293.52 552.50 l
	 292.65 528.47 l
	 290.03 528.47 l
	 280.42 528.47 l
	 279.76 545.94 l
	 276.70 545.94 l
	 277.36 532.84 l
	 278.89 526.28 l
	 289.81 526.28 l
	 288.94 506.62 l
	 284.35 506.62 l
	 281.51 521.91 l
	 270.80 519.73 l
	 270.37 528.47 l
	 270.58 535.02 l
cp p3
/bg { 1.0000 0.3647 0.0000 } def
np
  292.43 519.73 m
	 309.91 519.73 l
	 308.16 500.07 l
	 297.89 500.07 l
	 291.12 504.44 l
cp p3
/bg { 1.0000 0.4549 0.0000 } def
np
  312.97 552.50 m
	 332.41 552.50 l
	 331.97 497.88 l
	 308.16 500.07 l
	 309.91 519.73 l
cp p3
/bg { 1.0000 0.5451 0.0000 } def
np
  332.41 552.50 m
	 353.60 552.50 l
	 356.00 517.54 l
	 360.81 517.54 l
	 363.00 495.70 l
	 331.97 497.88 l
	 332.19 524.10 l
cp p3
/bg { 1.0000 0.6353 0.0000 } def
np
  245.02 510.99 m
	 245.90 513.17 l
	 261.19 510.99 l
	 264.90 493.51 l
	 248.52 493.51 l
cp p3
/bg { 1.0000 0.7255 0.0000 } def
np
  248.52 493.51 m
	 264.90 493.51 l
	 265.34 484.77 l
	 250.49 484.77 l
cp p3
/bg { 1.0000 0.8196 0.0000 } def
np
  250.49 484.77 m
	 255.95 484.77 l
	 261.41 458.56 l
	 257.26 456.37 l
	 257.26 458.56 l
	 257.48 460.74 l
	 257.91 465.11 l
	 257.91 467.30 l
	 257.48 469.48 l
	 255.73 471.67 l
	 253.11 471.67 l
cp p3
/bg { 1.0000 0.9098 0.0000 } def
np
  301.17 436.71 m
	 299.42 465.11 l
	 331.76 467.30 l
	 331.54 438.90 l
cp p3
/bg { 1.0000 1.0000 0.0000 } def
np
  294.62 497.88 m
	 331.76 495.70 l
	 331.76 467.30 l
	 299.42 465.11 l
cp p3
/bg { 0.9098 1.0000 0.0000 } def
np
  277.79 467.30 m
	 299.42 465.11 l
	 301.17 436.71 l
	 292.43 434.53 l
cp p3
/bg { 0.8196 1.0000 0.0000 } def
np
  261.19 510.99 m
	 285.88 506.62 l
	 286.10 506.62 l
	 294.62 497.88 l
	 299.42 465.11 l
	 277.79 467.30 l
	 276.05 469.48 l
	 268.84 484.77 l
	 265.34 484.77 l
	 264.90 493.51 l
cp p3
/bg { 0.7255 1.0000 0.0000 } def
np
  257.69 456.37 m
	 261.19 456.37 l
	 267.53 430.16 l
	 262.50 430.16 l
	 262.06 432.34 l
	 260.75 432.34 l
cp p3
/bg { 0.6353 1.0000 0.0000 } def
np
  262.94 427.97 m
	 269.49 427.97 l
	 276.70 430.16 l
	 277.14 425.79 l
	 293.30 430.16 l
	 306.63 386.46 l
	 272.99 377.72 l
	 262.94 425.79 l
cp p3
/bg { 0.5451 1.0000 0.0000 } def
np
  294.18 432.34 m
	 311.22 434.53 l
	 328.26 436.71 l
	 343.77 438.90 l
	 348.36 397.39 l
	 345.96 397.39 l
	 312.75 386.46 l
	 311.87 388.65 l
	 309.47 388.65 l
cp p3
/bg { 0.4549 1.0000 0.0000 } def
np
  315.81 334.03 m
	 315.81 342.77 l
	 316.46 353.69 l
	 317.34 360.25 l
	 318.43 368.99 l
	 317.12 377.72 l
	 314.28 384.28 l
	 312.75 386.46 l
	 341.80 395.20 l
	 349.45 395.20 l
	 350.76 384.28 l
	 351.42 382.09 l
	 375.45 377.72 l
	 372.83 366.80 l
	 371.30 344.95 l
	 371.08 334.03 l
cp p3
/bg { 0.3647 1.0000 0.0000 } def
np
  211.16 532.84 m
	 210.94 552.50 l
	 233.23 552.50 l
	 236.94 532.84 l
cp p3
/bg { 0.2745 1.0000 0.0000 } def
np
  211.38 480.40 m
	 210.94 532.84 l
	 226.02 532.84 l
	 235.63 484.77 l
	 230.60 482.59 l
	 220.34 482.59 l
cp p3
/bg { 0.1804 1.0000 0.0000 } def
np
  226.02 532.84 m
	 233.44 532.84 l
	 243.06 484.77 l
	 235.63 484.77 l
cp p3
/bg { 0.0902 1.0000 0.0000 } def
np
  243.06 484.77 m
	 233.44 532.84 l
	 237.81 532.84 l
	 243.06 508.81 l
	 246.12 484.77 l
cp p3
/bg { 0.0000 1.0000 0.0000 } def
np
  211.16 462.93 m
	 224.92 465.11 l
	 231.48 417.05 l
	 211.16 414.86 l
cp p3
/bg { 0.0000 1.0000 0.0902 } def
np
  229.51 432.34 m
	 249.39 436.71 l
	 260.32 419.23 l
	 231.48 417.05 l
cp p3
/bg { 0.0000 1.0000 0.1804 } def
np
  211.16 414.86 m
	 231.48 417.05 l
	 233.01 401.76 l
	 211.16 399.57 l
cp p3
/bg { 0.0000 1.0000 0.2745 } def
np
  231.48 417.05 m
	 260.32 419.23 l
	 264.25 403.94 l
	 233.01 401.76 l
cp p3
/bg { 0.0000 1.0000 0.3647 } def
np
  211.16 399.57 m
	 233.01 401.76 l
	 235.63 384.28 l
	 210.94 379.91 l
cp p3
/bg { 0.0000 1.0000 0.4549 } def
np
  233.01 401.76 m
	 264.25 403.94 l
	 269.71 379.91 l
	 255.95 377.72 l
	 255.07 382.09 l
	 252.45 384.28 l
	 247.86 386.46 l
	 246.12 390.83 l
	 234.76 388.65 l
cp p3
/bg { 0.0000 1.0000 0.5451 } def
np
  255.29 375.54 m
	 270.15 377.72 l
	 273.64 362.43 l
	 254.42 362.43 l
	 253.11 371.17 l
cp p3
/bg { 0.0000 1.0000 0.6353 } def
np
  210.94 379.91 m
	 230.60 382.09 l
	 230.82 375.54 l
	 234.54 373.36 l
	 235.85 375.54 l
	 235.85 371.17 l
	 210.94 371.17 l
cp p3
/bg { 0.0000 1.0000 0.7255 } def
np
  210.94 371.17 m
	 235.85 371.17 l
	 237.81 360.25 l
	 210.72 358.06 l
cp p3
/bg { 0.0000 1.0000 0.8196 } def
np
  210.72 358.06 m
	 237.81 360.25 l
	 241.75 334.03 l
	 211.16 334.03 l
cp p3
/bg { 0.0000 1.0000 0.9098 } def
np
  241.75 334.03 m
	 237.81 360.25 l
	 238.47 360.25 l
	 254.42 362.43 l
	 273.64 362.43 l
	 279.10 334.03 l
cp p3
/bg { 0.0000 1.0000 1.0000 } def
np
  272.99 377.72 m
	 278.45 377.72 l
	 280.85 362.43 l
	 281.07 358.06 l
	 277.14 358.06 l
cp p3
/bg { 0.0000 0.9098 1.0000 } def
np
  278.45 377.72 m
	 306.63 386.46 l
	 307.51 386.46 l
	 313.19 377.72 l
	 314.93 371.17 l
	 314.50 360.25 l
	 282.60 355.88 l
	 281.07 358.06 l
	 280.85 362.43 l
cp p3
/bg { 0.0000 0.8196 1.0000 } def
np
  286.75 334.03 m
	 282.60 355.88 l
	 314.50 360.25 l
	 313.40 349.32 l
	 312.09 344.95 l
	 311.44 334.03 l
cp p3
/bg { 0.0000 0.7255 1.0000 } def
np
  282.38 334.03 m
	 279.98 342.77 l
	 278.23 353.69 l
	 279.98 355.88 l
	 282.60 347.14 l
	 285.44 334.03 l
cp p3
/bg { 0.0000 0.6353 1.0000 } def
np
  343.77 438.90 m
	 357.75 438.90 l
	 361.47 412.68 l
	 348.80 410.49 l
	 350.76 399.57 l
	 348.36 397.39 l
cp p3
/bg { 0.0000 0.5451 1.0000 } def
np
  357.75 438.90 m
	 366.27 441.08 l
	 370.42 412.68 l
	 361.47 412.68 l
cp p3
/bg { 0.0000 0.4549 1.0000 } def
np
  366.27 441.08 m
	 383.75 441.08 l
	 389.43 441.08 l
	 394.46 441.08 l
	 388.99 432.34 l
	 390.30 427.97 l
	 398.61 425.79 l
	 390.96 414.86 l
	 370.42 412.68 l
cp p3
/bg { 0.0000 0.3647 1.0000 } def
np
  406.47 436.71 m
	 415.43 436.71 l
	 420.02 434.53 l
	 424.60 436.71 l
	 424.60 414.86 l
	 394.24 412.68 l
cp p3
/bg { 0.0000 0.2745 1.0000 } def
np
  394.24 412.68 m
	 424.60 414.86 l
	 425.48 390.83 l
	 382.44 393.02 l
	 387.90 401.76 l
cp p3
/bg { 0.0000 0.1804 1.0000 } def
np
  382.44 393.02 m
	 425.48 390.83 l
	 425.70 358.06 l
	 381.78 360.25 l
	 381.78 384.28 l
	 379.82 386.46 l
cp p3
/bg { 0.0000 0.0902 1.0000 } def
np
  386.37 334.03 m
	 386.59 344.95 l
	 388.99 351.51 l
	 390.96 360.25 l
	 425.70 358.06 l
	 425.26 349.32 l
	 425.70 334.03 l
cp p3
/bg { 0.0000 0.0000 1.0000 } def
np
  349.45 395.20 m
	 352.29 397.39 l
	 353.82 393.02 l
	 356.66 390.83 l
	 357.32 384.28 l
	 350.76 384.28 l
cp p3
/bg { 0.0902 0.0000 1.0000 } def
np
  356.66 390.83 m
	 368.24 388.65 l
	 371.52 390.83 l
	 375.01 399.57 l
	 384.41 401.76 l
	 379.82 390.83 l
	 375.23 379.91 l
	 357.32 384.28 l
cp p3
/bg { 0.1804 0.0000 1.0000 } def
np
  371.52 412.68 m
	 390.96 414.86 l
	 387.68 403.94 l
	 383.09 403.94 l
	 382.66 406.13 l
	 376.98 406.13 l
	 376.76 410.49 l
	 372.39 410.49 l
cp p3
/bg { 0.2745 0.0000 1.0000 } def
np
  333.07 495.70 m
	 335.25 497.88 l
	 336.56 497.88 l
	 348.36 495.70 l
	 348.14 493.51 l
	 348.80 482.59 l
	 333.28 480.40 l
cp p3
/bg { 0.3647 0.0000 1.0000 } def
np
  333.28 480.40 m
	 348.80 482.59 l
	 348.36 467.30 l
	 333.50 467.30 l
cp p3
/bg { 0.4549 0.0000 1.0000 } def
np
  348.36 495.70 m
	 361.90 495.70 l
	 361.90 443.26 l
	 348.36 441.08 l
	 348.36 467.30 l
	 348.80 482.59 l
	 348.14 493.51 l
cp p3
/bg { 0.5451 0.0000 1.0000 } def
np
  361.90 495.70 m
	 367.80 493.51 l
	 367.58 486.96 l
	 372.17 486.96 l
	 371.52 443.26 l
	 361.90 443.26 l
cp p3
/bg { 0.6353 0.0000 1.0000 } def
np
  371.52 443.26 m
	 371.95 467.30 l
	 386.37 467.30 l
	 386.37 447.63 l
	 381.78 447.63 l
	 381.35 445.45 l
	 375.23 445.45 l
	 373.70 443.26 l
cp p3
/bg { 0.7255 0.0000 1.0000 } def
np
  387.25 493.51 m
	 409.75 493.51 l
	 410.40 469.48 l
	 386.59 467.30 l
	 386.37 486.96 l
cp p3
/bg { 0.8196 0.0000 1.0000 } def
np
  386.59 467.30 m
	 410.40 469.48 l
	 413.46 452.00 l
	 404.50 452.00 l
	 403.85 445.45 l
	 388.56 445.45 l
	 386.37 447.63 l
	 386.37 467.30 l
cp p3
/bg { 0.9098 0.0000 1.0000 } def
np
  420.23 445.45 m
	 417.39 454.19 l
	 416.08 469.48 l
	 415.43 482.59 l
	 413.46 484.77 l
	 413.24 491.33 l
	 424.60 491.33 l
	 424.60 447.63 l
cp p3
/bg { 1.0000 0.0000 1.0000 } def
np
  353.60 552.50 m
	 366.05 552.50 l
	 367.58 517.54 l
	 355.79 517.54 l
cp p3
/bg { 1.0000 0.0000 0.9098 } def
np
  363.00 517.54 m
	 367.58 517.54 l
	 366.49 543.76 l
	 375.45 541.58 l
	 381.78 495.70 l
	 364.96 497.88 l
cp p3
/bg { 1.0000 0.0000 0.8196 } def
np
  366.05 552.50 m
	 377.41 552.50 l
	 378.07 548.13 l
	 378.29 543.76 l
	 383.09 543.76 l
	 387.03 532.84 l
	 376.98 530.65 l
	 375.45 541.58 l
	 366.49 543.76 l
cp p3
/bg { 1.0000 0.0000 0.7255 } def
np
  377.41 552.50 m
	 411.93 552.50 l
	 413.46 535.02 l
	 387.03 532.84 l
	 383.09 543.76 l
	 378.29 543.76 l
	 378.07 548.13 l
cp p3
/bg { 1.0000 0.0000 0.6353 } def
np
  413.46 535.02 m
	 413.46 515.36 l
	 411.50 515.36 l
	 382.44 510.99 l
	 380.47 532.84 l
	 387.03 532.84 l
cp p3
/bg { 1.0000 0.0000 0.5451 } def
np
  382.44 510.99 m
	 398.17 513.17 l
	 411.50 515.36 l
	 413.46 515.36 l
	 411.06 493.51 l
	 382.66 495.70 l
cp p3
/bg { 1.0000 0.0000 0.4549 } def
np
  413.24 552.50 m
	 424.82 552.50 l
	 424.82 537.21 l
	 415.21 537.21 l
cp p3
/bg { 1.0000 0.0000 0.3647 } def
np
  415.21 537.21 m
	 424.82 537.21 l
	 424.82 504.44 l
	 413.46 504.44 l
	 413.46 515.36 l
cp p3
/bg { 1.0000 0.0000 0.2745 } def
np
  413.46 504.44 m
	 424.82 504.44 l
	 424.60 491.33 l
	 413.24 491.33 l
	 411.71 497.88 l
cp p3
/bg { 1.0000 0.0000 0.1804 } def
np
  379.60 386.46 m
	 380.69 384.28 l
	 381.78 384.28 l
	 381.78 360.25 l
	 374.14 360.25 l
	 375.45 373.36 l
cp p3
/bg { 1.0000 0.0000 0.0902 } def
np
  241.31 530.65 m
	 270.80 535.02 l
	 270.37 528.47 l
	 264.90 524.10 l
	 243.93 517.54 l
	 242.84 524.10 l
cp p3
ep
%%Trailer
%%Pages: 1
%%EOF
