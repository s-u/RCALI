%!PS-Adobe-3.0 EPSF-3.0
%%DocumentNeededResources: font Helvetica
%%+ font Helvetica-Bold
%%+ font Helvetica-Oblique
%%+ font Helvetica-BoldOblique
%%+ font Symbol
%%Title: R Graphics Output
%%Creator: R Software
%%Pages: (atend)
%%BoundingBox: 156 322 439 520
%%EndComments
%%BeginProlog
/bp  { gs gs } def
% begin .ps.prolog
/gs  { gsave } def
/gr  { grestore } def
/ep  { showpage gr gr } def
/m   { moveto } def
/l   { lineto } def
/np  { newpath } def
/cp  { closepath } def
/f   { fill } def
/o   { stroke } def
/c   { newpath 0 360 arc } def
/r   { 3 index 3 index moveto 1 index 4 -1 roll
       lineto exch 1 index lineto lineto closepath } def
/p1  { stroke } def
/p2  { gsave bg setrgbcolor fill grestore newpath } def
/p3  { gsave bg setrgbcolor fill grestore stroke } def
/t   { 6 -2 roll moveto gsave rotate
       ps mul neg 0 2 1 roll rmoveto
       1 index stringwidth pop
       mul neg 0 rmoveto show grestore } def
/cl  { grestore gsave newpath 3 index 3 index moveto 1 index
       4 -1 roll lineto  exch 1 index lineto lineto
       closepath clip newpath } def
/rgb { setrgbcolor } def
/s   { scalefont setfont } def
/R   { /Font1 findfont } def
/B   { /Font2 findfont } def
/I   { /Font3 findfont } def
/BI  { /Font4 findfont } def
/S   { /Font5 findfont } def
1 setlinecap 1 setlinejoin
% end   .ps.prolog
%%IncludeResource: font Helvetica
/Helvetica findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font1 exch definefont pop
%%IncludeResource: font Helvetica-Bold
/Helvetica-Bold findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font2 exch definefont pop
%%IncludeResource: font Helvetica-Oblique
/Helvetica-Oblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font3 exch definefont pop
%%IncludeResource: font Helvetica-BoldOblique
/Helvetica-BoldOblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font4 exch definefont pop
%%IncludeResource: font Symbol
/Symbol findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  currentdict
  end
/Font5 exch definefont pop
%%EndProlog
%%Page: 1 1
bp
200.55 351.97 437.93 518.72 cl
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
273.89 417.09 m
364.58 417.09 l
o
np
364.58 417.09 m
369.87 511.17 l
o
np
369.87 511.17 m
268.60 511.17 l
o
np
268.60 511.17 m
273.89 417.09 l
o
np
244.93 358.15 m
273.89 417.09 l
o
np
268.60 511.17 m
229.59 512.54 l
o
np
229.59 512.54 m
244.93 358.15 l
o
np
393.54 358.15 m
408.88 512.54 l
o
np
408.88 512.54 m
369.87 511.17 l
o
np
364.58 417.09 m
393.54 358.15 l
o
np
244.93 358.15 m
393.54 358.15 l
o
np
408.88 512.54 m
229.59 512.54 l
o
155.91 321.73 439.37 520.16 cl
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
277.96 358.15 m
277.37 351.32 l
o
/ps 12 def R 12 s
276.77 339.98 (-1) 0.50 0.00 0.00 t
np
319.24 358.15 m
319.24 351.32 l
o
319.24 339.98 (0) 0.50 0.00 0.00 t
np
360.52 358.15 m
361.11 351.32 l
o
361.71 339.98 (1) 0.50 0.00 0.00 t
np
254.17 376.94 m
250.57 373.51 l
o
247.01 365.80 (-1) 0.50 0.00 0.00 t
np
262.92 394.75 m
259.77 391.71 l
o
256.65 384.39 (0) 0.50 0.00 0.00 t
np
269.59 408.34 m
266.79 405.61 l
o
264.01 398.59 (1) 0.50 0.00 0.00 t
np
242.56 382.03 m
236.32 379.46 l
o
229.82 372.48 (0.05) 0.50 0.00 0.00 t
np
239.68 411.01 m
233.14 408.95 l
o
226.32 402.50 (0.10) 0.50 0.00 0.00 t
np
236.58 442.26 m
229.71 440.80 l
o
222.53 434.96 (0.15) 0.50 0.00 0.00 t
np
233.22 476.05 m
225.99 475.29 l
o
218.42 470.19 (0.20) 0.50 0.00 0.00 t
200.55 351.97 437.93 518.72 cl
/bg { 0.7451 0.7451 0.7451 } def
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
  306.25 420.59 m
	 308.61 420.88 l
	 308.73 420.77 l
	 306.39 420.55 l
cp p3
np
  308.61 420.88 m
	 310.97 421.13 l
	 311.06 420.96 l
	 308.73 420.77 l
cp p3
np
  310.97 421.13 m
	 313.33 421.33 l
	 313.40 421.11 l
	 311.06 420.96 l
cp p3
np
  313.33 421.33 m
	 315.69 421.47 l
	 315.73 421.21 l
	 313.40 421.11 l
cp p3
np
  315.69 421.47 m
	 318.06 421.54 l
	 318.07 421.27 l
	 315.73 421.21 l
cp p3
np
  318.06 421.54 m
	 320.42 421.54 l
	 320.41 421.27 l
	 318.07 421.27 l
cp p3
np
  320.42 421.54 m
	 322.78 421.47 l
	 322.74 421.21 l
	 320.41 421.27 l
cp p3
np
  322.78 421.47 m
	 325.15 421.33 l
	 325.08 421.11 l
	 322.74 421.21 l
cp p3
np
  325.15 421.33 m
	 327.51 421.13 l
	 327.42 420.96 l
	 325.08 421.11 l
cp p3
np
  327.51 421.13 m
	 329.87 420.88 l
	 329.75 420.77 l
	 327.42 420.96 l
cp p3
np
  329.87 420.88 m
	 332.23 420.59 l
	 332.08 420.55 l
	 329.75 420.77 l
cp p3
np
  332.23 420.59 m
	 334.58 420.27 l
	 334.41 420.30 l
	 332.08 420.55 l
cp p3
np
  334.58 420.27 m
	 336.94 419.92 l
	 336.74 420.03 l
	 334.41 420.30 l
cp p3
np
  336.94 419.92 m
	 339.29 419.56 l
	 339.07 419.75 l
	 336.74 420.03 l
cp p3
np
  339.29 419.56 m
	 341.64 419.20 l
	 341.39 419.46 l
	 339.07 419.75 l
cp p3
np
  341.64 419.20 m
	 343.98 418.84 l
	 343.72 419.18 l
	 341.39 419.46 l
cp p3
np
  343.98 418.84 m
	 346.33 418.49 l
	 346.04 418.89 l
	 343.72 419.18 l
cp p3
np
  346.33 418.49 m
	 348.67 418.16 l
	 348.36 418.62 l
	 346.04 418.89 l
cp p3
np
  348.67 418.16 m
	 351.01 417.84 l
	 350.68 418.36 l
	 348.36 418.62 l
cp p3
np
  351.01 417.84 m
	 353.35 417.54 l
	 353.00 418.11 l
	 350.68 418.36 l
cp p3
np
  353.35 417.54 m
	 355.70 417.26 l
	 355.32 417.88 l
	 353.00 418.11 l
cp p3
np
  355.70 417.26 m
	 358.03 417.00 l
	 357.63 417.66 l
	 355.32 417.88 l
cp p3
np
  358.03 417.00 m
	 360.37 416.76 l
	 359.95 417.45 l
	 357.63 417.66 l
cp p3
np
  360.37 416.76 m
	 362.71 416.54 l
	 362.27 417.26 l
	 359.95 417.45 l
cp p3
np
  362.71 416.54 m
	 365.05 416.33 l
	 364.58 417.09 l
	 362.27 417.26 l
cp p3
np
  301.54 419.92 m
	 303.89 420.27 l
	 304.06 420.30 l
	 301.73 420.03 l
cp p3
np
  273.42 416.33 m
	 275.76 416.54 l
	 276.21 417.26 l
	 273.89 417.09 l
cp p3
np
  275.76 416.54 m
	 278.10 416.76 l
	 278.52 417.45 l
	 276.21 417.26 l
cp p3
np
  278.10 416.76 m
	 280.44 417.00 l
	 280.84 417.66 l
	 278.52 417.45 l
cp p3
np
  280.44 417.00 m
	 282.78 417.26 l
	 283.16 417.88 l
	 280.84 417.66 l
cp p3
np
  282.78 417.26 m
	 285.12 417.54 l
	 285.48 418.11 l
	 283.16 417.88 l
cp p3
np
  285.12 417.54 m
	 287.46 417.84 l
	 287.80 418.36 l
	 285.48 418.11 l
cp p3
np
  287.46 417.84 m
	 289.80 418.16 l
	 290.11 418.62 l
	 287.80 418.36 l
cp p3
np
  289.80 418.16 m
	 292.15 418.49 l
	 292.44 418.89 l
	 290.11 418.62 l
cp p3
np
  292.15 418.49 m
	 294.49 418.84 l
	 294.76 419.18 l
	 292.44 418.89 l
cp p3
np
  294.49 418.84 m
	 296.84 419.20 l
	 297.08 419.46 l
	 294.76 419.18 l
cp p3
np
  296.84 419.20 m
	 299.19 419.56 l
	 299.41 419.75 l
	 297.08 419.46 l
cp p3
np
  299.19 419.56 m
	 301.54 419.92 l
	 301.73 420.03 l
	 299.41 419.75 l
cp p3
np
  303.89 420.27 m
	 306.25 420.59 l
	 306.39 420.55 l
	 304.06 420.30 l
cp p3
np
  363.17 415.81 m
	 365.53 415.58 l
	 365.05 416.33 l
	 362.71 416.54 l
cp p3
np
  303.71 420.43 m
	 306.10 420.85 l
	 306.25 420.59 l
	 303.89 420.27 l
cp p3
np
  306.10 420.85 m
	 308.48 421.24 l
	 308.61 420.88 l
	 306.25 420.59 l
cp p3
np
  308.48 421.24 m
	 310.87 421.57 l
	 310.97 421.13 l
	 308.61 420.88 l
cp p3
np
  310.87 421.57 m
	 313.26 421.84 l
	 313.33 421.33 l
	 310.97 421.13 l
cp p3
np
  313.26 421.84 m
	 315.65 422.02 l
	 315.69 421.47 l
	 313.33 421.33 l
cp p3
np
  315.65 422.02 m
	 318.04 422.11 l
	 318.06 421.54 l
	 315.69 421.47 l
cp p3
np
  318.04 422.11 m
	 320.43 422.11 l
	 320.42 421.54 l
	 318.06 421.54 l
cp p3
np
  320.43 422.11 m
	 322.83 422.02 l
	 322.78 421.47 l
	 320.42 421.54 l
cp p3
np
  322.83 422.02 m
	 325.22 421.84 l
	 325.15 421.33 l
	 322.78 421.47 l
cp p3
np
  325.22 421.84 m
	 327.61 421.57 l
	 327.51 421.13 l
	 325.15 421.33 l
cp p3
np
  327.61 421.57 m
	 330.00 421.24 l
	 329.87 420.88 l
	 327.51 421.13 l
cp p3
np
  330.00 421.24 m
	 332.38 420.85 l
	 332.23 420.59 l
	 329.87 420.88 l
cp p3
np
  332.38 420.85 m
	 334.76 420.43 l
	 334.58 420.27 l
	 332.23 420.59 l
cp p3
np
  334.76 420.43 m
	 337.14 419.98 l
	 336.94 419.92 l
	 334.58 420.27 l
cp p3
np
  337.14 419.98 m
	 339.51 419.51 l
	 339.29 419.56 l
	 336.94 419.92 l
cp p3
np
  339.51 419.51 m
	 341.89 419.05 l
	 341.64 419.20 l
	 339.29 419.56 l
cp p3
np
  341.89 419.05 m
	 344.26 418.60 l
	 343.98 418.84 l
	 341.64 419.20 l
cp p3
np
  344.26 418.60 m
	 346.63 418.16 l
	 346.33 418.49 l
	 343.98 418.84 l
cp p3
np
  346.63 418.16 m
	 348.99 417.75 l
	 348.67 418.16 l
	 346.33 418.49 l
cp p3
np
  348.99 417.75 m
	 351.36 417.36 l
	 351.01 417.84 l
	 348.67 418.16 l
cp p3
np
  351.36 417.36 m
	 353.72 417.00 l
	 353.35 417.54 l
	 351.01 417.84 l
cp p3
np
  353.72 417.00 m
	 356.08 416.66 l
	 355.70 417.26 l
	 353.35 417.54 l
cp p3
np
  356.08 416.66 m
	 358.45 416.35 l
	 358.03 417.00 l
	 355.70 417.26 l
cp p3
np
  358.45 416.35 m
	 360.81 416.07 l
	 360.37 416.76 l
	 358.03 417.00 l
cp p3
np
  360.81 416.07 m
	 363.17 415.81 l
	 362.71 416.54 l
	 360.37 416.76 l
cp p3
np
  294.22 418.60 m
	 296.59 419.05 l
	 296.84 419.20 l
	 294.49 418.84 l
cp p3
np
  296.59 419.05 m
	 298.96 419.51 l
	 299.19 419.56 l
	 296.84 419.20 l
cp p3
np
  298.96 419.51 m
	 301.34 419.98 l
	 301.54 419.92 l
	 299.19 419.56 l
cp p3
np
  301.34 419.98 m
	 303.71 420.43 l
	 303.89 420.27 l
	 301.54 419.92 l
cp p3
np
  272.95 415.58 m
	 275.31 415.81 l
	 275.76 416.54 l
	 273.42 416.33 l
cp p3
np
  275.31 415.81 m
	 277.67 416.07 l
	 278.10 416.76 l
	 275.76 416.54 l
cp p3
np
  277.67 416.07 m
	 280.03 416.35 l
	 280.44 417.00 l
	 278.10 416.76 l
cp p3
np
  280.03 416.35 m
	 282.39 416.66 l
	 282.78 417.26 l
	 280.44 417.00 l
cp p3
np
  282.39 416.66 m
	 284.76 417.00 l
	 285.12 417.54 l
	 282.78 417.26 l
cp p3
np
  284.76 417.00 m
	 287.12 417.36 l
	 287.46 417.84 l
	 285.12 417.54 l
cp p3
np
  287.12 417.36 m
	 289.48 417.75 l
	 289.80 418.16 l
	 287.46 417.84 l
cp p3
np
  289.48 417.75 m
	 291.85 418.16 l
	 292.15 418.49 l
	 289.80 418.16 l
cp p3
np
  291.85 418.16 m
	 294.22 418.60 l
	 294.49 418.84 l
	 292.15 418.49 l
cp p3
np
  356.48 416.09 m
	 358.87 415.72 l
	 358.45 416.35 l
	 356.08 416.66 l
cp p3
np
  358.87 415.72 m
	 361.25 415.39 l
	 360.81 416.07 l
	 358.45 416.35 l
cp p3
np
  361.25 415.39 m
	 363.63 415.09 l
	 363.17 415.81 l
	 360.81 416.07 l
cp p3
np
  363.63 415.09 m
	 366.02 414.82 l
	 365.53 415.58 l
	 363.17 415.81 l
cp p3
np
  301.12 420.24 m
	 303.53 420.84 l
	 303.71 420.43 l
	 301.34 419.98 l
cp p3
np
  303.53 420.84 m
	 305.94 421.40 l
	 306.10 420.85 l
	 303.71 420.43 l
cp p3
np
  305.94 421.40 m
	 308.35 421.92 l
	 308.48 421.24 l
	 306.10 420.85 l
cp p3
np
  308.35 421.92 m
	 310.76 422.37 l
	 310.87 421.57 l
	 308.48 421.24 l
cp p3
np
  310.76 422.37 m
	 313.18 422.73 l
	 313.26 421.84 l
	 310.87 421.57 l
cp p3
np
  313.18 422.73 m
	 315.60 422.99 l
	 315.65 422.02 l
	 313.26 421.84 l
cp p3
np
  315.60 422.99 m
	 318.03 423.12 l
	 318.04 422.11 l
	 315.65 422.02 l
cp p3
np
  318.03 423.12 m
	 320.45 423.12 l
	 320.43 422.11 l
	 318.04 422.11 l
cp p3
np
  320.45 423.12 m
	 322.87 422.99 l
	 322.83 422.02 l
	 320.43 422.11 l
cp p3
np
  322.87 422.99 m
	 325.29 422.73 l
	 325.22 421.84 l
	 322.83 422.02 l
cp p3
np
  325.29 422.73 m
	 327.71 422.37 l
	 327.61 421.57 l
	 325.22 421.84 l
cp p3
np
  327.71 422.37 m
	 330.13 421.92 l
	 330.00 421.24 l
	 327.61 421.57 l
cp p3
np
  330.13 421.92 m
	 332.54 421.40 l
	 332.38 420.85 l
	 330.00 421.24 l
cp p3
np
  332.54 421.40 m
	 334.95 420.84 l
	 334.76 420.43 l
	 332.38 420.85 l
cp p3
np
  334.95 420.84 m
	 337.35 420.24 l
	 337.14 419.98 l
	 334.76 420.43 l
cp p3
np
  337.35 420.24 m
	 339.75 419.64 l
	 339.51 419.51 l
	 337.14 419.98 l
cp p3
np
  339.75 419.64 m
	 342.15 419.05 l
	 341.89 419.05 l
	 339.51 419.51 l
cp p3
np
  342.15 419.05 m
	 344.54 418.47 l
	 344.26 418.60 l
	 341.89 419.05 l
cp p3
np
  344.54 418.47 m
	 346.93 417.93 l
	 346.63 418.16 l
	 344.26 418.60 l
cp p3
np
  346.93 417.93 m
	 349.32 417.41 l
	 348.99 417.75 l
	 346.63 418.16 l
cp p3
np
  349.32 417.41 m
	 351.71 416.93 l
	 351.36 417.36 l
	 348.99 417.75 l
cp p3
np
  351.71 416.93 m
	 354.10 416.49 l
	 353.72 417.00 l
	 351.36 417.36 l
cp p3
np
  354.10 416.49 m
	 356.48 416.09 l
	 356.08 416.66 l
	 353.72 417.00 l
cp p3
np
  291.54 417.93 m
	 293.93 418.47 l
	 294.22 418.60 l
	 291.85 418.16 l
cp p3
np
  293.93 418.47 m
	 296.33 419.05 l
	 296.59 419.05 l
	 294.22 418.60 l
cp p3
np
  296.33 419.05 m
	 298.72 419.64 l
	 298.96 419.51 l
	 296.59 419.05 l
cp p3
np
  298.72 419.64 m
	 301.12 420.24 l
	 301.34 419.98 l
	 298.96 419.51 l
cp p3
np
  279.61 415.72 m
	 281.99 416.09 l
	 282.39 416.66 l
	 280.03 416.35 l
cp p3
np
  272.46 414.82 m
	 274.84 415.09 l
	 275.31 415.81 l
	 272.95 415.58 l
cp p3
np
  274.84 415.09 m
	 277.23 415.39 l
	 277.67 416.07 l
	 275.31 415.81 l
cp p3
np
  277.23 415.39 m
	 279.61 415.72 l
	 280.03 416.35 l
	 277.67 416.07 l
cp p3
np
  289.15 417.41 m
	 291.54 417.93 l
	 291.85 418.16 l
	 289.48 417.75 l
cp p3
np
  281.99 416.09 m
	 284.38 416.49 l
	 284.76 417.00 l
	 282.39 416.66 l
cp p3
np
  284.38 416.49 m
	 286.77 416.93 l
	 287.12 417.36 l
	 284.76 417.00 l
cp p3
np
  286.77 416.93 m
	 289.15 417.41 l
	 289.48 417.75 l
	 287.12 417.36 l
cp p3
np
  364.11 414.38 m
	 366.52 414.06 l
	 366.02 414.82 l
	 363.63 415.09 l
cp p3
np
  354.48 416.04 m
	 356.89 415.55 l
	 356.48 416.09 l
	 354.10 416.49 l
cp p3
np
  356.89 415.55 m
	 359.30 415.12 l
	 358.87 415.72 l
	 356.48 416.09 l
cp p3
np
  359.30 415.12 m
	 361.71 414.73 l
	 361.25 415.39 l
	 358.87 415.72 l
cp p3
np
  361.71 414.73 m
	 364.11 414.38 l
	 363.63 415.09 l
	 361.25 415.39 l
cp p3
np
  296.06 419.23 m
	 298.48 420.00 l
	 298.72 419.64 l
	 296.33 419.05 l
cp p3
np
  298.48 420.00 m
	 300.90 420.79 l
	 301.12 420.24 l
	 298.72 419.64 l
cp p3
np
  300.90 420.79 m
	 303.33 421.58 l
	 303.53 420.84 l
	 301.12 420.24 l
cp p3
np
  303.33 421.58 m
	 305.76 422.34 l
	 305.94 421.40 l
	 303.53 420.84 l
cp p3
np
  305.76 422.34 m
	 308.20 423.05 l
	 308.35 421.92 l
	 305.94 421.40 l
cp p3
np
  308.20 423.05 m
	 310.65 423.66 l
	 310.76 422.37 l
	 308.35 421.92 l
cp p3
np
  310.65 423.66 m
	 313.10 424.13 l
	 313.18 422.73 l
	 310.76 422.37 l
cp p3
np
  313.10 424.13 m
	 315.55 424.46 l
	 315.60 422.99 l
	 313.18 422.73 l
cp p3
np
  315.55 424.46 m
	 318.01 424.63 l
	 318.03 423.12 l
	 315.60 422.99 l
cp p3
np
  318.01 424.63 m
	 320.47 424.63 l
	 320.45 423.12 l
	 318.03 423.12 l
cp p3
np
  320.47 424.63 m
	 322.92 424.46 l
	 322.87 422.99 l
	 320.45 423.12 l
cp p3
np
  322.92 424.46 m
	 325.38 424.13 l
	 325.29 422.73 l
	 322.87 422.99 l
cp p3
np
  325.38 424.13 m
	 327.83 423.66 l
	 327.71 422.37 l
	 325.29 422.73 l
cp p3
np
  327.83 423.66 m
	 330.27 423.05 l
	 330.13 421.92 l
	 327.71 422.37 l
cp p3
np
  330.27 423.05 m
	 332.71 422.34 l
	 332.54 421.40 l
	 330.13 421.92 l
cp p3
np
  332.71 422.34 m
	 335.15 421.58 l
	 334.95 420.84 l
	 332.54 421.40 l
cp p3
np
  335.15 421.58 m
	 337.58 420.79 l
	 337.35 420.24 l
	 334.95 420.84 l
cp p3
np
  337.58 420.79 m
	 340.00 420.00 l
	 339.75 419.64 l
	 337.35 420.24 l
cp p3
np
  340.00 420.00 m
	 342.42 419.23 l
	 342.15 419.05 l
	 339.75 419.64 l
cp p3
np
  342.42 419.23 m
	 344.84 418.49 l
	 344.54 418.47 l
	 342.15 419.05 l
cp p3
np
  344.84 418.49 m
	 347.25 417.80 l
	 346.93 417.93 l
	 344.54 418.47 l
cp p3
np
  347.25 417.80 m
	 349.66 417.16 l
	 349.32 417.41 l
	 346.93 417.93 l
cp p3
np
  349.66 417.16 m
	 352.07 416.57 l
	 351.71 416.93 l
	 349.32 417.41 l
cp p3
np
  352.07 416.57 m
	 354.48 416.04 l
	 354.10 416.49 l
	 351.71 416.93 l
cp p3
np
  288.81 417.16 m
	 291.22 417.80 l
	 291.54 417.93 l
	 289.15 417.41 l
cp p3
np
  291.22 417.80 m
	 293.64 418.49 l
	 293.93 418.47 l
	 291.54 417.93 l
cp p3
np
  293.64 418.49 m
	 296.06 419.23 l
	 296.33 419.05 l
	 293.93 418.47 l
cp p3
np
  274.36 414.38 m
	 276.77 414.73 l
	 277.23 415.39 l
	 274.84 415.09 l
cp p3
np
  276.77 414.73 m
	 279.18 415.12 l
	 279.61 415.72 l
	 277.23 415.39 l
cp p3
np
  279.18 415.12 m
	 281.59 415.55 l
	 281.99 416.09 l
	 279.61 415.72 l
cp p3
np
  271.96 414.06 m
	 274.36 414.38 l
	 274.84 415.09 l
	 272.46 414.82 l
cp p3
np
  283.99 416.04 m
	 286.40 416.57 l
	 286.77 416.93 l
	 284.38 416.49 l
cp p3
np
  286.40 416.57 m
	 288.81 417.16 l
	 289.15 417.41 l
	 286.77 416.93 l
cp p3
np
  281.59 415.55 m
	 283.99 416.04 l
	 284.38 416.49 l
	 281.99 416.09 l
cp p3
np
  364.60 413.67 m
	 367.03 413.30 l
	 366.52 414.06 l
	 364.11 414.38 l
cp p3
np
  359.74 414.53 m
	 362.17 414.07 l
	 361.71 414.73 l
	 359.30 415.12 l
cp p3
np
  362.17 414.07 m
	 364.60 413.67 l
	 364.11 414.38 l
	 361.71 414.73 l
cp p3
np
  352.45 416.29 m
	 354.88 415.64 l
	 354.48 416.04 l
	 352.07 416.57 l
cp p3
np
  354.88 415.64 m
	 357.31 415.05 l
	 356.89 415.55 l
	 354.48 416.04 l
cp p3
np
  357.31 415.05 m
	 359.74 414.53 l
	 359.30 415.12 l
	 356.89 415.55 l
cp p3
np
  293.33 418.69 m
	 295.77 419.64 l
	 296.06 419.23 l
	 293.64 418.49 l
cp p3
np
  295.77 419.64 m
	 298.21 420.64 l
	 298.48 420.00 l
	 296.06 419.23 l
cp p3
np
  298.21 420.64 m
	 300.66 421.69 l
	 300.90 420.79 l
	 298.48 420.00 l
cp p3
np
  300.66 421.69 m
	 303.12 422.74 l
	 303.33 421.58 l
	 300.90 420.79 l
cp p3
np
  303.12 422.74 m
	 305.58 423.72 l
	 305.76 422.34 l
	 303.33 421.58 l
cp p3
np
  305.58 423.72 m
	 308.05 424.60 l
	 308.20 423.05 l
	 305.76 422.34 l
cp p3
np
  308.05 424.60 m
	 310.53 425.35 l
	 310.65 423.66 l
	 308.20 423.05 l
cp p3
np
  310.53 425.35 m
	 313.01 425.93 l
	 313.10 424.13 l
	 310.65 423.66 l
cp p3
np
  313.01 425.93 m
	 315.50 426.34 l
	 315.55 424.46 l
	 313.10 424.13 l
cp p3
np
  315.50 426.34 m
	 317.99 426.55 l
	 318.01 424.63 l
	 315.55 424.46 l
cp p3
np
  317.99 426.55 m
	 320.48 426.55 l
	 320.47 424.63 l
	 318.01 424.63 l
cp p3
np
  320.48 426.55 m
	 322.97 426.34 l
	 322.92 424.46 l
	 320.47 424.63 l
cp p3
np
  322.97 426.34 m
	 325.46 425.93 l
	 325.38 424.13 l
	 322.92 424.46 l
cp p3
np
  325.46 425.93 m
	 327.94 425.35 l
	 327.83 423.66 l
	 325.38 424.13 l
cp p3
np
  327.94 425.35 m
	 330.42 424.60 l
	 330.27 423.05 l
	 327.83 423.66 l
cp p3
np
  330.42 424.60 m
	 332.89 423.72 l
	 332.71 422.34 l
	 330.27 423.05 l
cp p3
np
  332.89 423.72 m
	 335.36 422.74 l
	 335.15 421.58 l
	 332.71 422.34 l
cp p3
np
  335.36 422.74 m
	 337.81 421.69 l
	 337.58 420.79 l
	 335.15 421.58 l
cp p3
np
  337.81 421.69 m
	 340.26 420.64 l
	 340.00 420.00 l
	 337.58 420.79 l
cp p3
np
  340.26 420.64 m
	 342.71 419.64 l
	 342.42 419.23 l
	 340.00 420.00 l
cp p3
np
  342.71 419.64 m
	 345.15 418.69 l
	 344.84 418.49 l
	 342.42 419.23 l
cp p3
np
  345.15 418.69 m
	 347.58 417.81 l
	 347.25 417.80 l
	 344.84 418.49 l
cp p3
np
  347.58 417.81 m
	 350.02 417.01 l
	 349.66 417.16 l
	 347.25 417.80 l
cp p3
np
  350.02 417.01 m
	 352.45 416.29 l
	 352.07 416.57 l
	 349.66 417.16 l
cp p3
np
  283.60 415.64 m
	 286.03 416.29 l
	 286.40 416.57 l
	 283.99 416.04 l
cp p3
np
  286.03 416.29 m
	 288.46 417.01 l
	 288.81 417.16 l
	 286.40 416.57 l
cp p3
np
  288.46 417.01 m
	 290.89 417.81 l
	 291.22 417.80 l
	 288.81 417.16 l
cp p3
np
  290.89 417.81 m
	 293.33 418.69 l
	 293.64 418.49 l
	 291.22 417.80 l
cp p3
np
  271.44 413.30 m
	 273.87 413.67 l
	 274.36 414.38 l
	 271.96 414.06 l
cp p3
np
  273.87 413.67 m
	 276.30 414.07 l
	 276.77 414.73 l
	 274.36 414.38 l
cp p3
np
  276.30 414.07 m
	 278.73 414.53 l
	 279.18 415.12 l
	 276.77 414.73 l
cp p3
np
  278.73 414.53 m
	 281.16 415.05 l
	 281.59 415.55 l
	 279.18 415.12 l
cp p3
np
  281.16 415.05 m
	 283.60 415.64 l
	 283.99 416.04 l
	 281.59 415.55 l
cp p3
np
  360.20 413.98 m
	 362.65 413.44 l
	 362.17 414.07 l
	 359.74 414.53 l
cp p3
np
  362.65 413.44 m
	 365.10 412.96 l
	 364.60 413.67 l
	 362.17 414.07 l
cp p3
np
  365.10 412.96 m
	 367.56 412.54 l
	 367.03 413.30 l
	 364.60 413.67 l
cp p3
np
  357.74 414.59 m
	 360.20 413.98 l
	 359.74 414.53 l
	 357.31 415.05 l
cp p3
np
  347.93 417.99 m
	 350.38 416.98 l
	 350.02 417.01 l
	 347.58 417.81 l
cp p3
np
  350.38 416.98 m
	 352.84 416.09 l
	 352.45 416.29 l
	 350.02 417.01 l
cp p3
np
  352.84 416.09 m
	 355.29 415.29 l
	 354.88 415.64 l
	 352.45 416.29 l
cp p3
np
  355.29 415.29 m
	 357.74 414.59 l
	 357.31 415.05 l
	 354.88 415.64 l
cp p3
np
  290.55 417.99 m
	 293.01 419.10 l
	 293.33 418.69 l
	 290.89 417.81 l
cp p3
np
  293.01 419.10 m
	 295.47 420.33 l
	 295.77 419.64 l
	 293.33 418.69 l
cp p3
np
  295.47 420.33 m
	 297.94 421.65 l
	 298.21 420.64 l
	 295.77 419.64 l
cp p3
np
  297.94 421.65 m
	 300.41 422.97 l
	 300.66 421.69 l
	 298.21 420.64 l
cp p3
np
  300.41 422.97 m
	 302.90 424.25 l
	 303.12 422.74 l
	 300.66 421.69 l
cp p3
np
  302.90 424.25 m
	 305.39 425.44 l
	 305.58 423.72 l
	 303.12 422.74 l
cp p3
np
  305.39 425.44 m
	 307.89 426.51 l
	 308.05 424.60 l
	 305.58 423.72 l
cp p3
np
  307.89 426.51 m
	 310.40 427.43 l
	 310.53 425.35 l
	 308.05 424.60 l
cp p3
np
  310.40 427.43 m
	 312.92 428.15 l
	 313.01 425.93 l
	 310.53 425.35 l
cp p3
np
  312.92 428.15 m
	 315.45 428.64 l
	 315.50 426.34 l
	 313.01 425.93 l
cp p3
np
  315.45 428.64 m
	 317.97 428.90 l
	 317.99 426.55 l
	 315.50 426.34 l
cp p3
np
  317.97 428.90 m
	 320.50 428.90 l
	 320.48 426.55 l
	 317.99 426.55 l
cp p3
np
  320.50 428.90 m
	 323.03 428.64 l
	 322.97 426.34 l
	 320.48 426.55 l
cp p3
np
  323.03 428.64 m
	 325.55 428.15 l
	 325.46 425.93 l
	 322.97 426.34 l
cp p3
np
  325.55 428.15 m
	 328.07 427.43 l
	 327.94 425.35 l
	 325.46 425.93 l
cp p3
np
  328.07 427.43 m
	 330.58 426.51 l
	 330.42 424.60 l
	 327.94 425.35 l
cp p3
np
  330.58 426.51 m
	 333.09 425.44 l
	 332.89 423.72 l
	 330.42 424.60 l
cp p3
np
  333.09 425.44 m
	 335.58 424.25 l
	 335.36 422.74 l
	 332.89 423.72 l
cp p3
np
  335.58 424.25 m
	 338.06 422.97 l
	 337.81 421.69 l
	 335.36 422.74 l
cp p3
np
  338.06 422.97 m
	 340.54 421.65 l
	 340.26 420.64 l
	 337.81 421.69 l
cp p3
np
  340.54 421.65 m
	 343.01 420.33 l
	 342.71 419.64 l
	 340.26 420.64 l
cp p3
np
  343.01 420.33 m
	 345.47 419.10 l
	 345.15 418.69 l
	 342.71 419.64 l
cp p3
np
  345.47 419.10 m
	 347.93 417.99 l
	 347.58 417.81 l
	 345.15 418.69 l
cp p3
np
  280.73 414.59 m
	 283.19 415.29 l
	 283.60 415.64 l
	 281.16 415.05 l
cp p3
np
  283.19 415.29 m
	 285.64 416.09 l
	 286.03 416.29 l
	 283.60 415.64 l
cp p3
np
  285.64 416.09 m
	 288.09 416.98 l
	 288.46 417.01 l
	 286.03 416.29 l
cp p3
np
  288.09 416.98 m
	 290.55 417.99 l
	 290.89 417.81 l
	 288.46 417.01 l
cp p3
np
  278.28 413.98 m
	 280.73 414.59 l
	 281.16 415.05 l
	 278.73 414.53 l
cp p3
np
  270.92 412.54 m
	 273.37 412.96 l
	 273.87 413.67 l
	 271.44 413.30 l
cp p3
np
  273.37 412.96 m
	 275.83 413.44 l
	 276.30 414.07 l
	 273.87 413.67 l
cp p3
np
  275.83 413.44 m
	 278.28 413.98 l
	 278.73 414.53 l
	 276.30 414.07 l
cp p3
np
  355.71 415.02 m
	 358.19 414.17 l
	 357.74 414.59 l
	 355.29 415.29 l
cp p3
np
  358.19 414.17 m
	 360.66 413.44 l
	 360.20 413.98 l
	 357.74 414.59 l
cp p3
np
  360.66 413.44 m
	 363.14 412.81 l
	 362.65 413.44 l
	 360.20 413.98 l
cp p3
np
  363.14 412.81 m
	 365.62 412.26 l
	 365.10 412.96 l
	 362.65 413.44 l
cp p3
np
  365.62 412.26 m
	 368.09 411.78 l
	 367.56 412.54 l
	 365.10 412.96 l
cp p3
np
  345.81 419.79 m
	 348.29 418.36 l
	 347.93 417.99 l
	 345.47 419.10 l
cp p3
np
  348.29 418.36 m
	 350.76 417.09 l
	 350.38 416.98 l
	 347.93 417.99 l
cp p3
np
  350.76 417.09 m
	 353.24 415.98 l
	 352.84 416.09 l
	 350.38 416.98 l
cp p3
np
  353.24 415.98 m
	 355.71 415.02 l
	 355.29 415.29 l
	 352.84 416.09 l
cp p3
np
  285.24 415.98 m
	 287.71 417.09 l
	 288.09 416.98 l
	 285.64 416.09 l
cp p3
np
  287.71 417.09 m
	 290.19 418.36 l
	 290.55 417.99 l
	 288.09 416.98 l
cp p3
np
  290.19 418.36 m
	 292.67 419.79 l
	 293.01 419.10 l
	 290.55 417.99 l
cp p3
np
  292.67 419.79 m
	 295.15 421.35 l
	 295.47 420.33 l
	 293.01 419.10 l
cp p3
np
  295.15 421.35 m
	 297.65 422.94 l
	 297.94 421.65 l
	 295.47 420.33 l
cp p3
np
  297.65 422.94 m
	 300.15 424.52 l
	 300.41 422.97 l
	 297.94 421.65 l
cp p3
np
  300.15 424.52 m
	 302.66 426.06 l
	 302.90 424.25 l
	 300.41 422.97 l
cp p3
np
  302.66 426.06 m
	 305.19 427.50 l
	 305.39 425.44 l
	 302.90 424.25 l
cp p3
np
  305.19 427.50 m
	 307.72 428.80 l
	 307.89 426.51 l
	 305.39 425.44 l
cp p3
np
  307.72 428.80 m
	 310.27 429.91 l
	 310.40 427.43 l
	 307.89 426.51 l
cp p3
np
  310.27 429.91 m
	 312.83 430.78 l
	 312.92 428.15 l
	 310.40 427.43 l
cp p3
np
  312.83 430.78 m
	 315.39 431.39 l
	 315.45 428.64 l
	 312.92 428.15 l
cp p3
np
  315.39 431.39 m
	 317.95 431.70 l
	 317.97 428.90 l
	 315.45 428.64 l
cp p3
np
  317.95 431.70 m
	 320.52 431.70 l
	 320.50 428.90 l
	 317.97 428.90 l
cp p3
np
  320.52 431.70 m
	 323.09 431.39 l
	 323.03 428.64 l
	 320.50 428.90 l
cp p3
np
  323.09 431.39 m
	 325.65 430.78 l
	 325.55 428.15 l
	 323.03 428.64 l
cp p3
np
  325.65 430.78 m
	 328.21 429.91 l
	 328.07 427.43 l
	 325.55 428.15 l
cp p3
np
  328.21 429.91 m
	 330.75 428.80 l
	 330.58 426.51 l
	 328.07 427.43 l
cp p3
np
  330.75 428.80 m
	 333.29 427.50 l
	 333.09 425.44 l
	 330.58 426.51 l
cp p3
np
  333.29 427.50 m
	 335.81 426.06 l
	 335.58 424.25 l
	 333.09 425.44 l
cp p3
np
  335.81 426.06 m
	 338.33 424.52 l
	 338.06 422.97 l
	 335.58 424.25 l
cp p3
np
  338.33 424.52 m
	 340.83 422.94 l
	 340.54 421.65 l
	 338.06 422.97 l
cp p3
np
  340.83 422.94 m
	 343.32 421.35 l
	 343.01 420.33 l
	 340.54 421.65 l
cp p3
np
  343.32 421.35 m
	 345.81 419.79 l
	 345.47 419.10 l
	 343.01 420.33 l
cp p3
np
  277.81 413.44 m
	 280.29 414.17 l
	 280.73 414.59 l
	 278.28 413.98 l
cp p3
np
  280.29 414.17 m
	 282.76 415.02 l
	 283.19 415.29 l
	 280.73 414.59 l
cp p3
np
  282.76 415.02 m
	 285.24 415.98 l
	 285.64 416.09 l
	 283.19 415.29 l
cp p3
np
  272.86 412.26 m
	 275.34 412.81 l
	 275.83 413.44 l
	 273.37 412.96 l
cp p3
np
  275.34 412.81 m
	 277.81 413.44 l
	 278.28 413.98 l
	 275.83 413.44 l
cp p3
np
  270.38 411.78 m
	 272.86 412.26 l
	 273.37 412.96 l
	 270.92 412.54 l
cp p3
np
  356.15 414.81 m
	 358.65 413.80 l
	 358.19 414.17 l
	 355.71 415.02 l
cp p3
np
  351.16 417.36 m
	 353.65 415.99 l
	 353.24 415.98 l
	 350.76 417.09 l
cp p3
np
  353.65 415.99 m
	 356.15 414.81 l
	 355.71 415.02 l
	 353.24 415.98 l
cp p3
np
  366.14 411.56 m
	 368.64 411.01 l
	 368.09 411.78 l
	 365.62 412.26 l
cp p3
np
  358.65 413.80 m
	 361.14 412.94 l
	 360.66 413.44 l
	 358.19 414.17 l
cp p3
np
  361.14 412.94 m
	 363.64 412.20 l
	 363.14 412.81 l
	 360.66 413.44 l
cp p3
np
  363.64 412.20 m
	 366.14 411.56 l
	 365.62 412.26 l
	 363.14 412.81 l
cp p3
np
  343.65 422.56 m
	 346.16 420.72 l
	 345.81 419.79 l
	 343.32 421.35 l
cp p3
np
  346.16 420.72 m
	 348.66 418.95 l
	 348.29 418.36 l
	 345.81 419.79 l
cp p3
np
  348.66 418.95 m
	 351.16 417.36 l
	 350.76 417.09 l
	 348.29 418.36 l
cp p3
np
  282.33 414.81 m
	 284.82 415.99 l
	 285.24 415.98 l
	 282.76 415.02 l
cp p3
np
  284.82 415.99 m
	 287.32 417.36 l
	 287.71 417.09 l
	 285.24 415.98 l
cp p3
np
  287.32 417.36 m
	 289.81 418.95 l
	 290.19 418.36 l
	 287.71 417.09 l
cp p3
np
  289.81 418.95 m
	 292.31 420.72 l
	 292.67 419.79 l
	 290.19 418.36 l
cp p3
np
  292.31 420.72 m
	 294.82 422.56 l
	 295.15 421.35 l
	 292.67 419.79 l
cp p3
np
  294.82 422.56 m
	 297.34 424.45 l
	 297.65 422.94 l
	 295.15 421.35 l
cp p3
np
  297.34 424.45 m
	 299.87 426.34 l
	 300.15 424.52 l
	 297.65 422.94 l
cp p3
np
  299.87 426.34 m
	 302.42 428.18 l
	 302.66 426.06 l
	 300.15 424.52 l
cp p3
np
  302.42 428.18 m
	 304.97 429.91 l
	 305.19 427.50 l
	 302.66 426.06 l
cp p3
np
  304.97 429.91 m
	 307.55 431.47 l
	 307.72 428.80 l
	 305.19 427.50 l
cp p3
np
  307.55 431.47 m
	 310.13 432.80 l
	 310.27 429.91 l
	 307.72 428.80 l
cp p3
np
  310.13 432.80 m
	 312.72 433.86 l
	 312.83 430.78 l
	 310.27 429.91 l
cp p3
np
  312.72 433.86 m
	 315.33 434.60 l
	 315.39 431.39 l
	 312.83 430.78 l
cp p3
np
  315.33 434.60 m
	 317.93 434.97 l
	 317.95 431.70 l
	 315.39 431.39 l
cp p3
np
  317.93 434.97 m
	 320.54 434.97 l
	 320.52 431.70 l
	 317.95 431.70 l
cp p3
np
  320.54 434.97 m
	 323.15 434.60 l
	 323.09 431.39 l
	 320.52 431.70 l
cp p3
np
  323.15 434.60 m
	 325.75 433.86 l
	 325.65 430.78 l
	 323.09 431.39 l
cp p3
np
  325.75 433.86 m
	 328.35 432.80 l
	 328.21 429.91 l
	 325.65 430.78 l
cp p3
np
  328.35 432.80 m
	 330.93 431.47 l
	 330.75 428.80 l
	 328.21 429.91 l
cp p3
np
  330.93 431.47 m
	 333.50 429.91 l
	 333.29 427.50 l
	 330.75 428.80 l
cp p3
np
  333.50 429.91 m
	 336.06 428.18 l
	 335.81 426.06 l
	 333.29 427.50 l
cp p3
np
  336.06 428.18 m
	 338.60 426.34 l
	 338.33 424.52 l
	 335.81 426.06 l
cp p3
np
  338.60 426.34 m
	 341.14 424.45 l
	 340.83 422.94 l
	 338.33 424.52 l
cp p3
np
  341.14 424.45 m
	 343.65 422.56 l
	 343.32 421.35 l
	 340.83 422.94 l
cp p3
np
  272.33 411.56 m
	 274.83 412.20 l
	 275.34 412.81 l
	 272.86 412.26 l
cp p3
np
  274.83 412.20 m
	 277.33 412.94 l
	 277.81 413.44 l
	 275.34 412.81 l
cp p3
np
  277.33 412.94 m
	 279.83 413.80 l
	 280.29 414.17 l
	 277.81 413.44 l
cp p3
np
  279.83 413.80 m
	 282.33 414.81 l
	 282.76 415.02 l
	 280.29 414.17 l
cp p3
np
  269.83 411.01 m
	 272.33 411.56 l
	 272.86 412.26 l
	 270.38 411.78 l
cp p3
np
  351.57 417.79 m
	 354.09 416.10 l
	 353.65 415.99 l
	 351.16 417.36 l
cp p3
np
  354.09 416.10 m
	 356.60 414.67 l
	 356.15 414.81 l
	 353.65 415.99 l
cp p3
np
  356.60 414.67 m
	 359.12 413.47 l
	 358.65 413.80 l
	 356.15 414.81 l
cp p3
np
  349.06 419.73 m
	 351.57 417.79 l
	 351.16 417.36 l
	 348.66 418.95 l
cp p3
np
  361.64 412.45 m
	 364.16 411.59 l
	 363.64 412.20 l
	 361.14 412.94 l
cp p3
np
  364.16 411.59 m
	 366.68 410.86 l
	 366.14 411.56 l
	 363.64 412.20 l
cp p3
np
  366.68 410.86 m
	 369.21 410.24 l
	 368.64 411.01 l
	 366.14 411.56 l
cp p3
np
  359.12 413.47 m
	 361.64 412.45 l
	 361.14 412.94 l
	 358.65 413.80 l
cp p3
np
  338.89 428.41 m
	 341.45 426.18 l
	 341.14 424.45 l
	 338.60 426.34 l
cp p3
np
  341.45 426.18 m
	 344.00 423.96 l
	 343.65 422.56 l
	 341.14 424.45 l
cp p3
np
  344.00 423.96 m
	 346.53 421.79 l
	 346.16 420.72 l
	 343.65 422.56 l
cp p3
np
  346.53 421.79 m
	 349.06 419.73 l
	 348.66 418.95 l
	 346.16 420.72 l
cp p3
np
  279.36 413.47 m
	 281.88 414.67 l
	 282.33 414.81 l
	 279.83 413.80 l
cp p3
np
  281.88 414.67 m
	 284.39 416.10 l
	 284.82 415.99 l
	 282.33 414.81 l
cp p3
np
  284.39 416.10 m
	 286.90 417.79 l
	 287.32 417.36 l
	 284.82 415.99 l
cp p3
np
  286.90 417.79 m
	 289.42 419.73 l
	 289.81 418.95 l
	 287.32 417.36 l
cp p3
np
  289.42 419.73 m
	 291.94 421.79 l
	 292.31 420.72 l
	 289.81 418.95 l
cp p3
np
  291.94 421.79 m
	 294.48 423.96 l
	 294.82 422.56 l
	 292.31 420.72 l
cp p3
np
  294.48 423.96 m
	 297.02 426.18 l
	 297.34 424.45 l
	 294.82 422.56 l
cp p3
np
  297.02 426.18 m
	 299.58 428.41 l
	 299.87 426.34 l
	 297.34 424.45 l
cp p3
np
  299.58 428.41 m
	 302.16 430.59 l
	 302.42 428.18 l
	 299.87 426.34 l
cp p3
np
  302.16 430.59 m
	 304.75 432.65 l
	 304.97 429.91 l
	 302.42 428.18 l
cp p3
np
  304.75 432.65 m
	 307.36 434.52 l
	 307.55 431.47 l
	 304.97 429.91 l
cp p3
np
  307.36 434.52 m
	 309.98 436.13 l
	 310.13 432.80 l
	 307.55 431.47 l
cp p3
np
  309.98 436.13 m
	 312.61 437.41 l
	 312.72 433.86 l
	 310.13 432.80 l
cp p3
np
  312.61 437.41 m
	 315.26 438.30 l
	 315.33 434.60 l
	 312.72 433.86 l
cp p3
np
  315.26 438.30 m
	 317.91 438.76 l
	 317.93 434.97 l
	 315.33 434.60 l
cp p3
np
  317.91 438.76 m
	 320.56 438.76 l
	 320.54 434.97 l
	 317.93 434.97 l
cp p3
np
  320.56 438.76 m
	 323.22 438.30 l
	 323.15 434.60 l
	 320.54 434.97 l
cp p3
np
  323.22 438.30 m
	 325.86 437.41 l
	 325.75 433.86 l
	 323.15 434.60 l
cp p3
np
  325.86 437.41 m
	 328.50 436.13 l
	 328.35 432.80 l
	 325.75 433.86 l
cp p3
np
  328.50 436.13 m
	 331.12 434.52 l
	 330.93 431.47 l
	 328.35 432.80 l
cp p3
np
  331.12 434.52 m
	 333.73 432.65 l
	 333.50 429.91 l
	 330.93 431.47 l
cp p3
np
  333.73 432.65 m
	 336.32 430.59 l
	 336.06 428.18 l
	 333.50 429.91 l
cp p3
np
  336.32 430.59 m
	 338.89 428.41 l
	 338.60 426.34 l
	 336.06 428.18 l
cp p3
np
  269.27 410.24 m
	 271.79 410.86 l
	 272.33 411.56 l
	 269.83 411.01 l
cp p3
np
  271.79 410.86 m
	 274.32 411.59 l
	 274.83 412.20 l
	 272.33 411.56 l
cp p3
np
  274.32 411.59 m
	 276.84 412.45 l
	 277.33 412.94 l
	 274.83 412.20 l
cp p3
np
  276.84 412.45 m
	 279.36 413.47 l
	 279.83 413.80 l
	 277.33 412.94 l
cp p3
np
  346.92 422.99 m
	 349.46 420.60 l
	 349.06 419.73 l
	 346.53 421.79 l
cp p3
np
  349.46 420.60 m
	 352.00 418.37 l
	 351.57 417.79 l
	 349.06 419.73 l
cp p3
np
  352.00 418.37 m
	 354.53 416.33 l
	 354.09 416.10 l
	 351.57 417.79 l
cp p3
np
  354.53 416.33 m
	 357.07 414.61 l
	 356.60 414.67 l
	 354.09 416.10 l
cp p3
np
  357.07 414.61 m
	 359.60 413.17 l
	 359.12 413.47 l
	 356.60 414.67 l
cp p3
np
  359.60 413.17 m
	 362.14 411.98 l
	 361.64 412.45 l
	 359.12 413.47 l
cp p3
np
  362.14 411.98 m
	 364.69 410.99 l
	 364.16 411.59 l
	 361.64 412.45 l
cp p3
np
  364.69 410.99 m
	 367.23 410.15 l
	 366.68 410.86 l
	 364.16 411.59 l
cp p3
np
  367.23 410.15 m
	 369.78 409.45 l
	 369.21 410.24 l
	 366.68 410.86 l
cp p3
np
  336.59 433.27 m
	 339.20 430.70 l
	 338.89 428.41 l
	 336.32 430.59 l
cp p3
np
  339.20 430.70 m
	 341.78 428.09 l
	 341.45 426.18 l
	 338.89 428.41 l
cp p3
np
  341.78 428.09 m
	 344.36 425.51 l
	 344.00 423.96 l
	 341.45 426.18 l
cp p3
np
  344.36 425.51 m
	 346.92 422.99 l
	 346.53 421.79 l
	 344.00 423.96 l
cp p3
np
  271.24 410.15 m
	 273.79 410.99 l
	 274.32 411.59 l
	 271.79 410.86 l
cp p3
np
  273.79 410.99 m
	 276.33 411.98 l
	 276.84 412.45 l
	 274.32 411.59 l
cp p3
np
  276.33 411.98 m
	 278.87 413.17 l
	 279.36 413.47 l
	 276.84 412.45 l
cp p3
np
  278.87 413.17 m
	 281.41 414.61 l
	 281.88 414.67 l
	 279.36 413.47 l
cp p3
np
  281.41 414.61 m
	 283.94 416.33 l
	 284.39 416.10 l
	 281.88 414.67 l
cp p3
np
  283.94 416.33 m
	 286.48 418.37 l
	 286.90 417.79 l
	 284.39 416.10 l
cp p3
np
  286.48 418.37 m
	 289.01 420.60 l
	 289.42 419.73 l
	 286.90 417.79 l
cp p3
np
  289.01 420.60 m
	 291.56 422.99 l
	 291.94 421.79 l
	 289.42 419.73 l
cp p3
np
  291.56 422.99 m
	 294.12 425.51 l
	 294.48 423.96 l
	 291.94 421.79 l
cp p3
np
  294.12 425.51 m
	 296.69 428.09 l
	 297.02 426.18 l
	 294.48 423.96 l
cp p3
np
  296.69 428.09 m
	 299.28 430.70 l
	 299.58 428.41 l
	 297.02 426.18 l
cp p3
np
  299.28 430.70 m
	 301.89 433.27 l
	 302.16 430.59 l
	 299.58 428.41 l
cp p3
np
  301.89 433.27 m
	 304.51 435.71 l
	 304.75 432.65 l
	 302.16 430.59 l
cp p3
np
  304.51 435.71 m
	 307.16 437.94 l
	 307.36 434.52 l
	 304.75 432.65 l
cp p3
np
  307.16 437.94 m
	 309.82 439.88 l
	 309.98 436.13 l
	 307.36 434.52 l
cp p3
np
  309.82 439.88 m
	 312.50 441.43 l
	 312.61 437.41 l
	 309.98 436.13 l
cp p3
np
  312.50 441.43 m
	 315.19 442.52 l
	 315.26 438.30 l
	 312.61 437.41 l
cp p3
np
  315.19 442.52 m
	 317.89 443.07 l
	 317.91 438.76 l
	 315.26 438.30 l
cp p3
np
  317.89 443.07 m
	 320.59 443.07 l
	 320.56 438.76 l
	 317.91 438.76 l
cp p3
np
  320.59 443.07 m
	 323.29 442.52 l
	 323.22 438.30 l
	 320.56 438.76 l
cp p3
np
  323.29 442.52 m
	 325.98 441.43 l
	 325.86 437.41 l
	 323.22 438.30 l
cp p3
np
  325.98 441.43 m
	 328.66 439.88 l
	 328.50 436.13 l
	 325.86 437.41 l
cp p3
np
  328.66 439.88 m
	 331.32 437.94 l
	 331.12 434.52 l
	 328.50 436.13 l
cp p3
np
  331.32 437.94 m
	 333.96 435.71 l
	 333.73 432.65 l
	 331.12 434.52 l
cp p3
np
  333.96 435.71 m
	 336.59 433.27 l
	 336.32 430.59 l
	 333.73 432.65 l
cp p3
np
  268.69 409.45 m
	 271.24 410.15 l
	 271.79 410.86 l
	 269.27 410.24 l
cp p3
np
  334.21 439.07 m
	 336.87 436.18 l
	 336.59 433.27 l
	 333.96 435.71 l
cp p3
np
  339.51 433.18 m
	 342.13 430.15 l
	 341.78 428.09 l
	 339.20 430.70 l
cp p3
np
  342.13 430.15 m
	 344.73 427.16 l
	 344.36 425.51 l
	 341.78 428.09 l
cp p3
np
  344.73 427.16 m
	 347.31 424.27 l
	 346.92 422.99 l
	 344.36 425.51 l
cp p3
np
  347.31 424.27 m
	 349.88 421.54 l
	 349.46 420.60 l
	 346.92 422.99 l
cp p3
np
  349.88 421.54 m
	 352.44 418.99 l
	 352.00 418.37 l
	 349.46 420.60 l
cp p3
np
  352.44 418.99 m
	 354.99 416.66 l
	 354.53 416.33 l
	 352.00 418.37 l
cp p3
np
  354.99 416.66 m
	 357.54 414.60 l
	 357.07 414.61 l
	 354.53 416.33 l
cp p3
np
  357.54 414.60 m
	 360.10 412.91 l
	 359.60 413.17 l
	 357.07 414.61 l
cp p3
np
  360.10 412.91 m
	 362.66 411.52 l
	 362.14 411.98 l
	 359.60 413.17 l
cp p3
np
  362.66 411.52 m
	 365.23 410.38 l
	 364.69 410.99 l
	 362.14 411.98 l
cp p3
np
  365.23 410.38 m
	 367.80 409.43 l
	 367.23 410.15 l
	 364.69 410.99 l
cp p3
np
  367.80 409.43 m
	 370.37 408.64 l
	 369.78 409.45 l
	 367.23 410.15 l
cp p3
np
  336.87 436.18 m
	 339.51 433.18 l
	 339.20 430.70 l
	 336.59 433.27 l
cp p3
np
  268.10 408.64 m
	 270.68 409.43 l
	 271.24 410.15 l
	 268.69 409.45 l
cp p3
np
  270.68 409.43 m
	 273.25 410.38 l
	 273.79 410.99 l
	 271.24 410.15 l
cp p3
np
  273.25 410.38 m
	 275.81 411.52 l
	 276.33 411.98 l
	 273.79 410.99 l
cp p3
np
  275.81 411.52 m
	 278.37 412.91 l
	 278.87 413.17 l
	 276.33 411.98 l
cp p3
np
  278.37 412.91 m
	 280.93 414.60 l
	 281.41 414.61 l
	 278.87 413.17 l
cp p3
np
  280.93 414.60 m
	 283.48 416.66 l
	 283.94 416.33 l
	 281.41 414.61 l
cp p3
np
  283.48 416.66 m
	 286.03 418.99 l
	 286.48 418.37 l
	 283.94 416.33 l
cp p3
np
  286.03 418.99 m
	 288.59 421.54 l
	 289.01 420.60 l
	 286.48 418.37 l
cp p3
np
  288.59 421.54 m
	 291.16 424.27 l
	 291.56 422.99 l
	 289.01 420.60 l
cp p3
np
  291.16 424.27 m
	 293.75 427.16 l
	 294.12 425.51 l
	 291.56 422.99 l
cp p3
np
  293.75 427.16 m
	 296.35 430.15 l
	 296.69 428.09 l
	 294.12 425.51 l
cp p3
np
  296.35 430.15 m
	 298.97 433.18 l
	 299.28 430.70 l
	 296.69 428.09 l
cp p3
np
  298.97 433.18 m
	 301.60 436.18 l
	 301.89 433.27 l
	 299.28 430.70 l
cp p3
np
  301.60 436.18 m
	 304.27 439.07 l
	 304.51 435.71 l
	 301.89 433.27 l
cp p3
np
  304.27 439.07 m
	 306.95 441.73 l
	 307.16 437.94 l
	 304.51 435.71 l
cp p3
np
  306.95 441.73 m
	 309.65 444.06 l
	 309.82 439.88 l
	 307.16 437.94 l
cp p3
np
  309.65 444.06 m
	 312.38 445.95 l
	 312.50 441.43 l
	 309.82 439.88 l
cp p3
np
  312.38 445.95 m
	 315.11 447.28 l
	 315.19 442.52 l
	 312.50 441.43 l
cp p3
np
  315.11 447.28 m
	 317.86 447.96 l
	 317.89 443.07 l
	 315.19 442.52 l
cp p3
np
  317.86 447.96 m
	 320.61 447.96 l
	 320.59 443.07 l
	 317.89 443.07 l
cp p3
np
  320.61 447.96 m
	 323.36 447.28 l
	 323.29 442.52 l
	 320.59 443.07 l
cp p3
np
  323.36 447.28 m
	 326.10 445.95 l
	 325.98 441.43 l
	 323.29 442.52 l
cp p3
np
  326.10 445.95 m
	 328.82 444.06 l
	 328.66 439.88 l
	 325.98 441.43 l
cp p3
np
  328.82 444.06 m
	 331.53 441.73 l
	 331.32 437.94 l
	 328.66 439.88 l
cp p3
np
  331.53 441.73 m
	 334.21 439.07 l
	 333.96 435.71 l
	 331.32 437.94 l
cp p3
np
  326.23 450.97 m
	 329.00 448.67 l
	 328.82 444.06 l
	 326.10 445.95 l
cp p3
np
  329.00 448.67 m
	 331.75 445.86 l
	 331.53 441.73 l
	 328.82 444.06 l
cp p3
np
  331.75 445.86 m
	 334.47 442.68 l
	 334.21 439.07 l
	 331.53 441.73 l
cp p3
np
  334.47 442.68 m
	 337.16 439.28 l
	 336.87 436.18 l
	 334.21 439.07 l
cp p3
np
  337.16 439.28 m
	 339.84 435.78 l
	 339.51 433.18 l
	 336.87 436.18 l
cp p3
np
  339.84 435.78 m
	 342.48 432.28 l
	 342.13 430.15 l
	 339.51 433.18 l
cp p3
np
  342.48 432.28 m
	 345.11 428.86 l
	 344.73 427.16 l
	 342.13 430.15 l
cp p3
np
  345.11 428.86 m
	 347.72 425.58 l
	 347.31 424.27 l
	 344.73 427.16 l
cp p3
np
  347.72 425.58 m
	 350.31 422.49 l
	 349.88 421.54 l
	 347.31 424.27 l
cp p3
np
  350.31 422.49 m
	 352.89 419.61 l
	 352.44 418.99 l
	 349.88 421.54 l
cp p3
np
  352.89 419.61 m
	 355.47 416.99 l
	 354.99 416.66 l
	 352.44 418.99 l
cp p3
np
  355.47 416.99 m
	 358.04 414.63 l
	 357.54 414.60 l
	 354.99 416.66 l
cp p3
np
  358.04 414.63 m
	 360.61 412.66 l
	 360.10 412.91 l
	 357.54 414.60 l
cp p3
np
  360.61 412.66 m
	 363.19 411.06 l
	 362.66 411.52 l
	 360.10 412.91 l
cp p3
np
  363.19 411.06 m
	 365.78 409.76 l
	 365.23 410.38 l
	 362.66 411.52 l
cp p3
np
  365.78 409.76 m
	 368.38 408.69 l
	 367.80 409.43 l
	 365.23 410.38 l
cp p3
np
  368.38 408.69 m
	 370.98 407.80 l
	 370.37 408.64 l
	 367.80 409.43 l
cp p3
np
  298.64 435.78 m
	 301.31 439.28 l
	 301.60 436.18 l
	 298.97 433.18 l
cp p3
np
  267.50 407.80 m
	 270.10 408.69 l
	 270.68 409.43 l
	 268.10 408.64 l
cp p3
np
  270.10 408.69 m
	 272.69 409.76 l
	 273.25 410.38 l
	 270.68 409.43 l
cp p3
np
  272.69 409.76 m
	 275.28 411.06 l
	 275.81 411.52 l
	 273.25 410.38 l
cp p3
np
  275.28 411.06 m
	 277.86 412.66 l
	 278.37 412.91 l
	 275.81 411.52 l
cp p3
np
  277.86 412.66 m
	 280.44 414.63 l
	 280.93 414.60 l
	 278.37 412.91 l
cp p3
np
  280.44 414.63 m
	 283.01 416.99 l
	 283.48 416.66 l
	 280.93 414.60 l
cp p3
np
  283.01 416.99 m
	 285.58 419.61 l
	 286.03 418.99 l
	 283.48 416.66 l
cp p3
np
  285.58 419.61 m
	 288.16 422.49 l
	 288.59 421.54 l
	 286.03 418.99 l
cp p3
np
  288.16 422.49 m
	 290.76 425.58 l
	 291.16 424.27 l
	 288.59 421.54 l
cp p3
np
  290.76 425.58 m
	 293.37 428.86 l
	 293.75 427.16 l
	 291.16 424.27 l
cp p3
np
  293.37 428.86 m
	 295.99 432.28 l
	 296.35 430.15 l
	 293.75 427.16 l
cp p3
np
  295.99 432.28 m
	 298.64 435.78 l
	 298.97 433.18 l
	 296.35 430.15 l
cp p3
np
  309.48 448.67 m
	 312.25 450.97 l
	 312.38 445.95 l
	 309.65 444.06 l
cp p3
np
  301.31 439.28 m
	 304.01 442.68 l
	 304.27 439.07 l
	 301.60 436.18 l
cp p3
np
  304.01 442.68 m
	 306.73 445.86 l
	 306.95 441.73 l
	 304.27 439.07 l
cp p3
np
  306.73 445.86 m
	 309.48 448.67 l
	 309.65 444.06 l
	 306.95 441.73 l
cp p3
np
  320.64 453.46 m
	 323.44 452.61 l
	 323.36 447.28 l
	 320.61 447.96 l
cp p3
np
  312.25 450.97 m
	 315.03 452.61 l
	 315.11 447.28 l
	 312.38 445.95 l
cp p3
np
  315.03 452.61 m
	 317.84 453.46 l
	 317.86 447.96 l
	 315.11 447.28 l
cp p3
np
  317.84 453.46 m
	 320.64 453.46 l
	 320.61 447.96 l
	 317.86 447.96 l
cp p3
np
  323.44 452.61 m
	 326.23 450.97 l
	 326.10 445.95 l
	 323.36 447.28 l
cp p3
np
  368.97 407.91 m
	 371.59 406.94 l
	 370.98 407.80 l
	 368.38 408.69 l
cp p3
np
  323.53 458.54 m
	 326.37 456.50 l
	 326.23 450.97 l
	 323.44 452.61 l
cp p3
np
  326.37 456.50 m
	 329.19 453.67 l
	 329.00 448.67 l
	 326.23 450.97 l
cp p3
np
  329.19 453.67 m
	 331.98 450.26 l
	 331.75 445.86 l
	 329.00 448.67 l
cp p3
np
  331.98 450.26 m
	 334.74 446.48 l
	 334.47 442.68 l
	 331.75 445.86 l
cp p3
np
  334.74 446.48 m
	 337.47 442.49 l
	 337.16 439.28 l
	 334.47 442.68 l
cp p3
np
  337.47 442.49 m
	 340.17 438.44 l
	 339.84 435.78 l
	 337.16 439.28 l
cp p3
np
  340.17 438.44 m
	 342.85 434.43 l
	 342.48 432.28 l
	 339.84 435.78 l
cp p3
np
  342.85 434.43 m
	 345.50 430.55 l
	 345.11 428.86 l
	 342.48 432.28 l
cp p3
np
  345.50 430.55 m
	 348.13 426.86 l
	 347.72 425.58 l
	 345.11 428.86 l
cp p3
np
  348.13 426.86 m
	 350.75 423.40 l
	 350.31 422.49 l
	 347.72 425.58 l
cp p3
np
  350.75 423.40 m
	 353.36 420.20 l
	 352.89 419.61 l
	 350.31 422.49 l
cp p3
np
  353.36 420.20 m
	 355.95 417.28 l
	 355.47 416.99 l
	 352.89 419.61 l
cp p3
np
  355.95 417.28 m
	 358.55 414.67 l
	 358.04 414.63 l
	 355.47 416.99 l
cp p3
np
  358.55 414.67 m
	 361.14 412.40 l
	 360.61 412.66 l
	 358.04 414.63 l
cp p3
np
  361.14 412.40 m
	 363.74 410.57 l
	 363.19 411.06 l
	 360.61 412.66 l
cp p3
np
  363.74 410.57 m
	 366.35 409.11 l
	 365.78 409.76 l
	 363.19 411.06 l
cp p3
np
  366.35 409.11 m
	 368.97 407.91 l
	 368.38 408.69 l
	 365.78 409.76 l
cp p3
np
  292.98 430.55 m
	 295.63 434.43 l
	 295.99 432.28 l
	 293.37 428.86 l
cp p3
np
  295.63 434.43 m
	 298.31 438.44 l
	 298.64 435.78 l
	 295.99 432.28 l
cp p3
np
  298.31 438.44 m
	 301.01 442.49 l
	 301.31 439.28 l
	 298.64 435.78 l
cp p3
np
  266.88 406.94 m
	 269.51 407.91 l
	 270.10 408.69 l
	 267.50 407.80 l
cp p3
np
  269.51 407.91 m
	 272.13 409.11 l
	 272.69 409.76 l
	 270.10 408.69 l
cp p3
np
  272.13 409.11 m
	 274.74 410.57 l
	 275.28 411.06 l
	 272.69 409.76 l
cp p3
np
  274.74 410.57 m
	 277.34 412.40 l
	 277.86 412.66 l
	 275.28 411.06 l
cp p3
np
  277.34 412.40 m
	 279.93 414.67 l
	 280.44 414.63 l
	 277.86 412.66 l
cp p3
np
  279.93 414.67 m
	 282.52 417.28 l
	 283.01 416.99 l
	 280.44 414.63 l
cp p3
np
  282.52 417.28 m
	 285.12 420.20 l
	 285.58 419.61 l
	 283.01 416.99 l
cp p3
np
  285.12 420.20 m
	 287.72 423.40 l
	 288.16 422.49 l
	 285.58 419.61 l
cp p3
np
  287.72 423.40 m
	 290.34 426.86 l
	 290.76 425.58 l
	 288.16 422.49 l
cp p3
np
  290.34 426.86 m
	 292.98 430.55 l
	 293.37 428.86 l
	 290.76 425.58 l
cp p3
np
  303.74 446.48 m
	 306.50 450.26 l
	 306.73 445.86 l
	 304.01 442.68 l
cp p3
np
  306.50 450.26 m
	 309.29 453.67 l
	 309.48 448.67 l
	 306.73 445.86 l
cp p3
np
  309.29 453.67 m
	 312.11 456.50 l
	 312.25 450.97 l
	 309.48 448.67 l
cp p3
np
  301.01 442.49 m
	 303.74 446.48 l
	 304.01 442.68 l
	 301.31 439.28 l
cp p3
np
  314.95 458.54 m
	 317.81 459.62 l
	 317.84 453.46 l
	 315.03 452.61 l
cp p3
np
  317.81 459.62 m
	 320.67 459.62 l
	 320.64 453.46 l
	 317.84 453.46 l
cp p3
np
  320.67 459.62 m
	 323.53 458.54 l
	 323.44 452.61 l
	 320.64 453.46 l
cp p3
np
  312.11 456.50 m
	 314.95 458.54 l
	 315.03 452.61 l
	 312.25 450.97 l
cp p3
np
  364.30 410.04 m
	 366.93 408.41 l
	 366.35 409.11 l
	 363.74 410.57 l
cp p3
np
  366.93 408.41 m
	 369.57 407.09 l
	 368.97 407.91 l
	 366.35 409.11 l
cp p3
np
  369.57 407.09 m
	 372.22 406.03 l
	 371.59 406.94 l
	 368.97 407.91 l
cp p3
np
  320.70 466.47 m
	 323.62 465.09 l
	 323.53 458.54 l
	 320.67 459.62 l
cp p3
np
  323.62 465.09 m
	 326.51 462.51 l
	 326.37 456.50 l
	 323.53 458.54 l
cp p3
np
  326.51 462.51 m
	 329.38 459.00 l
	 329.19 453.67 l
	 326.37 456.50 l
cp p3
np
  329.38 459.00 m
	 332.22 454.86 l
	 331.98 450.26 l
	 329.19 453.67 l
cp p3
np
  332.22 454.86 m
	 335.01 450.36 l
	 334.74 446.48 l
	 331.98 450.26 l
cp p3
np
  335.01 450.36 m
	 337.78 445.71 l
	 337.47 442.49 l
	 334.74 446.48 l
cp p3
np
  337.78 445.71 m
	 340.51 441.05 l
	 340.17 438.44 l
	 337.47 442.49 l
cp p3
np
  340.51 441.05 m
	 343.22 436.51 l
	 342.85 434.43 l
	 340.17 438.44 l
cp p3
np
  343.22 436.51 m
	 345.90 432.15 l
	 345.50 430.55 l
	 342.85 434.43 l
cp p3
np
  345.90 432.15 m
	 348.56 428.04 l
	 348.13 426.86 l
	 345.50 430.55 l
cp p3
np
  348.56 428.04 m
	 351.20 424.21 l
	 350.75 423.40 l
	 348.13 426.86 l
cp p3
np
  351.20 424.21 m
	 353.83 420.69 l
	 353.36 420.20 l
	 350.75 423.40 l
cp p3
np
  353.83 420.69 m
	 356.45 417.49 l
	 355.95 417.28 l
	 353.36 420.20 l
cp p3
np
  356.45 417.49 m
	 359.06 414.62 l
	 358.55 414.67 l
	 355.95 417.28 l
cp p3
np
  359.06 414.62 m
	 361.68 412.10 l
	 361.14 412.40 l
	 358.55 414.67 l
cp p3
np
  361.68 412.10 m
	 364.30 410.04 l
	 363.74 410.57 l
	 361.14 412.40 l
cp p3
np
  289.92 428.04 m
	 292.58 432.15 l
	 292.98 430.55 l
	 290.34 426.86 l
cp p3
np
  292.58 432.15 m
	 295.26 436.51 l
	 295.63 434.43 l
	 292.98 430.55 l
cp p3
np
  295.26 436.51 m
	 297.96 441.05 l
	 298.31 438.44 l
	 295.63 434.43 l
cp p3
np
  297.96 441.05 m
	 300.70 445.71 l
	 301.01 442.49 l
	 298.31 438.44 l
cp p3
np
  266.25 406.03 m
	 268.90 407.09 l
	 269.51 407.91 l
	 266.88 406.94 l
cp p3
np
  268.90 407.09 m
	 271.55 408.41 l
	 272.13 409.11 l
	 269.51 407.91 l
cp p3
np
  271.55 408.41 m
	 274.18 410.04 l
	 274.74 410.57 l
	 272.13 409.11 l
cp p3
np
  274.18 410.04 m
	 276.80 412.10 l
	 277.34 412.40 l
	 274.74 410.57 l
cp p3
np
  276.80 412.10 m
	 279.41 414.62 l
	 279.93 414.67 l
	 277.34 412.40 l
cp p3
np
  279.41 414.62 m
	 282.03 417.49 l
	 282.52 417.28 l
	 279.93 414.67 l
cp p3
np
  282.03 417.49 m
	 284.65 420.69 l
	 285.12 420.20 l
	 282.52 417.28 l
cp p3
np
  284.65 420.69 m
	 287.28 424.21 l
	 287.72 423.40 l
	 285.12 420.20 l
cp p3
np
  287.28 424.21 m
	 289.92 428.04 l
	 290.34 426.86 l
	 287.72 423.40 l
cp p3
np
  300.70 445.71 m
	 303.46 450.36 l
	 303.74 446.48 l
	 301.01 442.49 l
cp p3
np
  303.46 450.36 m
	 306.26 454.86 l
	 306.50 450.26 l
	 303.74 446.48 l
cp p3
np
  306.26 454.86 m
	 309.09 459.00 l
	 309.29 453.67 l
	 306.50 450.26 l
cp p3
np
  309.09 459.00 m
	 311.96 462.51 l
	 312.11 456.50 l
	 309.29 453.67 l
cp p3
np
  311.96 462.51 m
	 314.86 465.09 l
	 314.95 458.54 l
	 312.11 456.50 l
cp p3
np
  314.86 465.09 m
	 317.78 466.47 l
	 317.81 459.62 l
	 314.95 458.54 l
cp p3
np
  317.78 466.47 m
	 320.70 466.47 l
	 320.67 459.62 l
	 317.81 459.62 l
cp p3
np
  370.19 406.22 m
	 372.87 405.06 l
	 372.22 406.03 l
	 369.57 407.09 l
cp p3
np
  362.22 411.74 m
	 364.87 409.45 l
	 364.30 410.04 l
	 361.68 412.10 l
cp p3
np
  364.87 409.45 m
	 367.52 407.65 l
	 366.93 408.41 l
	 364.30 410.04 l
cp p3
np
  367.52 407.65 m
	 370.19 406.22 l
	 369.57 407.09 l
	 366.93 408.41 l
cp p3
np
  314.76 472.26 m
	 317.74 474.07 l
	 317.78 466.47 l
	 314.86 465.09 l
cp p3
np
  317.74 474.07 m
	 320.73 474.07 l
	 320.70 466.47 l
	 317.78 466.47 l
cp p3
np
  320.73 474.07 m
	 323.71 472.26 l
	 323.62 465.09 l
	 320.70 466.47 l
cp p3
np
  323.71 472.26 m
	 326.67 468.92 l
	 326.51 462.51 l
	 323.62 465.09 l
cp p3
np
  326.67 468.92 m
	 329.58 464.53 l
	 329.38 459.00 l
	 326.51 462.51 l
cp p3
np
  329.58 464.53 m
	 332.46 459.50 l
	 332.22 454.86 l
	 329.38 459.00 l
cp p3
np
  332.46 459.50 m
	 335.30 454.18 l
	 335.01 450.36 l
	 332.22 454.86 l
cp p3
np
  335.30 454.18 m
	 338.10 448.79 l
	 337.78 445.71 l
	 335.01 450.36 l
cp p3
np
  338.10 448.79 m
	 340.86 443.49 l
	 340.51 441.05 l
	 337.78 445.71 l
cp p3
np
  340.86 443.49 m
	 343.59 438.40 l
	 343.22 436.51 l
	 340.51 441.05 l
cp p3
np
  343.59 438.40 m
	 346.30 433.57 l
	 345.90 432.15 l
	 343.22 436.51 l
cp p3
np
  346.30 433.57 m
	 348.99 429.05 l
	 348.56 428.04 l
	 345.90 432.15 l
cp p3
np
  348.99 429.05 m
	 351.65 424.86 l
	 351.20 424.21 l
	 348.56 428.04 l
cp p3
np
  351.65 424.86 m
	 354.31 421.03 l
	 353.83 420.69 l
	 351.20 424.21 l
cp p3
np
  354.31 421.03 m
	 356.95 417.56 l
	 356.45 417.49 l
	 353.83 420.69 l
cp p3
np
  356.95 417.56 m
	 359.59 414.46 l
	 359.06 414.62 l
	 356.45 417.49 l
cp p3
np
  359.59 414.46 m
	 362.22 411.74 l
	 361.68 412.10 l
	 359.06 414.62 l
cp p3
np
  286.82 424.86 m
	 289.49 429.05 l
	 289.92 428.04 l
	 287.28 424.21 l
cp p3
np
  289.49 429.05 m
	 292.17 433.57 l
	 292.58 432.15 l
	 289.92 428.04 l
cp p3
np
  292.17 433.57 m
	 294.88 438.40 l
	 295.26 436.51 l
	 292.58 432.15 l
cp p3
np
  294.88 438.40 m
	 297.61 443.49 l
	 297.96 441.05 l
	 295.26 436.51 l
cp p3
np
  297.61 443.49 m
	 300.38 448.79 l
	 300.70 445.71 l
	 297.96 441.05 l
cp p3
np
  265.61 405.06 m
	 268.29 406.22 l
	 268.90 407.09 l
	 266.25 406.03 l
cp p3
np
  268.29 406.22 m
	 270.95 407.65 l
	 271.55 408.41 l
	 268.90 407.09 l
cp p3
np
  270.95 407.65 m
	 273.61 409.45 l
	 274.18 410.04 l
	 271.55 408.41 l
cp p3
np
  273.61 409.45 m
	 276.25 411.74 l
	 276.80 412.10 l
	 274.18 410.04 l
cp p3
np
  276.25 411.74 m
	 278.89 414.46 l
	 279.41 414.62 l
	 276.80 412.10 l
cp p3
np
  278.89 414.46 m
	 281.53 417.56 l
	 282.03 417.49 l
	 279.41 414.62 l
cp p3
np
  281.53 417.56 m
	 284.17 421.03 l
	 284.65 420.69 l
	 282.03 417.49 l
cp p3
np
  284.17 421.03 m
	 286.82 424.86 l
	 287.28 424.21 l
	 284.65 420.69 l
cp p3
np
  308.89 464.53 m
	 311.81 468.92 l
	 311.96 462.51 l
	 309.09 459.00 l
cp p3
np
  300.38 448.79 m
	 303.18 454.18 l
	 303.46 450.36 l
	 300.70 445.71 l
cp p3
np
  303.18 454.18 m
	 306.01 459.50 l
	 306.26 454.86 l
	 303.46 450.36 l
cp p3
np
  306.01 459.50 m
	 308.89 464.53 l
	 309.09 459.00 l
	 306.26 454.86 l
cp p3
np
  311.81 468.92 m
	 314.76 472.26 l
	 314.86 465.09 l
	 311.96 462.51 l
cp p3
np
  360.12 414.15 m
	 362.78 411.24 l
	 362.22 411.74 l
	 359.59 414.46 l
cp p3
np
  365.44 408.76 m
	 368.13 406.81 l
	 367.52 407.65 l
	 364.87 409.45 l
cp p3
np
  368.13 406.81 m
	 370.82 405.27 l
	 370.19 406.22 l
	 367.52 407.65 l
cp p3
np
  370.82 405.27 m
	 373.52 404.04 l
	 372.87 405.06 l
	 370.19 406.22 l
cp p3
np
  362.78 411.24 m
	 365.44 408.76 l
	 364.87 409.45 l
	 362.22 411.74 l
cp p3
np
  311.65 475.58 m
	 314.66 479.98 l
	 314.76 472.26 l
	 311.81 468.92 l
cp p3
np
  314.66 479.98 m
	 317.71 482.48 l
	 317.74 474.07 l
	 314.76 472.26 l
cp p3
np
  317.71 482.48 m
	 320.77 482.48 l
	 320.73 474.07 l
	 317.74 474.07 l
cp p3
np
  320.77 482.48 m
	 323.81 479.98 l
	 323.71 472.26 l
	 320.73 474.07 l
cp p3
np
  323.81 479.98 m
	 326.82 475.58 l
	 326.67 468.92 l
	 323.71 472.26 l
cp p3
np
  326.82 475.58 m
	 329.79 470.04 l
	 329.58 464.53 l
	 326.67 468.92 l
cp p3
np
  329.79 470.04 m
	 332.71 463.95 l
	 332.46 459.50 l
	 329.58 464.53 l
cp p3
np
  332.71 463.95 m
	 335.58 457.71 l
	 335.30 454.18 l
	 332.46 459.50 l
cp p3
np
  335.58 457.71 m
	 338.42 451.55 l
	 338.10 448.79 l
	 335.30 454.18 l
cp p3
np
  338.42 451.55 m
	 341.21 445.61 l
	 340.86 443.49 l
	 338.10 448.79 l
cp p3
np
  341.21 445.61 m
	 343.97 439.98 l
	 343.59 438.40 l
	 340.86 443.49 l
cp p3
np
  343.97 439.98 m
	 346.71 434.70 l
	 346.30 433.57 l
	 343.59 438.40 l
cp p3
np
  346.71 434.70 m
	 349.42 429.79 l
	 348.99 429.05 l
	 346.30 433.57 l
cp p3
np
  349.42 429.79 m
	 352.11 425.28 l
	 351.65 424.86 l
	 348.99 429.05 l
cp p3
np
  352.11 425.28 m
	 354.79 421.17 l
	 354.31 421.03 l
	 351.65 424.86 l
cp p3
np
  354.79 421.17 m
	 357.45 417.46 l
	 356.95 417.56 l
	 354.31 421.03 l
cp p3
np
  357.45 417.46 m
	 360.12 414.15 l
	 359.59 414.46 l
	 356.95 417.56 l
cp p3
np
  281.02 417.46 m
	 283.69 421.17 l
	 284.17 421.03 l
	 281.53 417.56 l
cp p3
np
  283.69 421.17 m
	 286.37 425.28 l
	 286.82 424.86 l
	 284.17 421.03 l
cp p3
np
  286.37 425.28 m
	 289.06 429.79 l
	 289.49 429.05 l
	 286.82 424.86 l
cp p3
np
  289.06 429.79 m
	 291.77 434.70 l
	 292.17 433.57 l
	 289.49 429.05 l
cp p3
np
  291.77 434.70 m
	 294.50 439.98 l
	 294.88 438.40 l
	 292.17 433.57 l
cp p3
np
  294.50 439.98 m
	 297.27 445.61 l
	 297.61 443.49 l
	 294.88 438.40 l
cp p3
np
  297.27 445.61 m
	 300.06 451.55 l
	 300.38 448.79 l
	 297.61 443.49 l
cp p3
np
  264.95 404.04 m
	 267.66 405.27 l
	 268.29 406.22 l
	 265.61 405.06 l
cp p3
np
  267.66 405.27 m
	 270.35 406.81 l
	 270.95 407.65 l
	 268.29 406.22 l
cp p3
np
  270.35 406.81 m
	 273.03 408.76 l
	 273.61 409.45 l
	 270.95 407.65 l
cp p3
np
  273.03 408.76 m
	 275.70 411.24 l
	 276.25 411.74 l
	 273.61 409.45 l
cp p3
np
  275.70 411.24 m
	 278.36 414.15 l
	 278.89 414.46 l
	 276.25 411.74 l
cp p3
np
  278.36 414.15 m
	 281.02 417.46 l
	 281.53 417.56 l
	 278.89 414.46 l
cp p3
np
  302.89 457.71 m
	 305.76 463.95 l
	 306.01 459.50 l
	 303.18 454.18 l
cp p3
np
  305.76 463.95 m
	 308.68 470.04 l
	 308.89 464.53 l
	 306.01 459.50 l
cp p3
np
  308.68 470.04 m
	 311.65 475.58 l
	 311.81 468.92 l
	 308.89 464.53 l
cp p3
np
  300.06 451.55 m
	 302.89 457.71 l
	 303.18 454.18 l
	 300.38 448.79 l
cp p3
np
  355.27 421.05 m
	 357.96 417.13 l
	 357.45 417.46 l
	 354.79 421.17 l
cp p3
np
  357.96 417.13 m
	 360.65 413.64 l
	 360.12 414.15 l
	 357.45 417.46 l
cp p3
np
  360.65 413.64 m
	 363.34 410.58 l
	 362.78 411.24 l
	 360.12 414.15 l
cp p3
np
  363.34 410.58 m
	 366.03 407.95 l
	 365.44 408.76 l
	 362.78 411.24 l
cp p3
np
  366.03 407.95 m
	 368.74 405.87 l
	 368.13 406.81 l
	 365.44 408.76 l
cp p3
np
  368.74 405.87 m
	 371.46 404.24 l
	 370.82 405.27 l
	 368.13 406.81 l
cp p3
np
  371.46 404.24 m
	 374.19 402.94 l
	 373.52 404.04 l
	 370.82 405.27 l
cp p3
np
  308.48 475.13 m
	 311.49 482.12 l
	 311.65 475.58 l
	 308.68 470.04 l
cp p3
np
  311.49 482.12 m
	 314.56 488.07 l
	 314.66 479.98 l
	 311.65 475.58 l
cp p3
np
  314.56 488.07 m
	 317.67 491.72 l
	 317.71 482.48 l
	 314.66 479.98 l
cp p3
np
  317.67 491.72 m
	 320.80 491.72 l
	 320.77 482.48 l
	 317.71 482.48 l
cp p3
np
  320.80 491.72 m
	 323.92 488.07 l
	 323.81 479.98 l
	 320.77 482.48 l
cp p3
np
  323.92 488.07 m
	 326.99 482.12 l
	 326.82 475.58 l
	 323.81 479.98 l
cp p3
np
  326.99 482.12 m
	 330.00 475.13 l
	 329.79 470.04 l
	 326.82 475.58 l
cp p3
np
  330.00 475.13 m
	 332.96 467.86 l
	 332.71 463.95 l
	 329.79 470.04 l
cp p3
np
  332.96 467.86 m
	 335.87 460.68 l
	 335.58 457.71 l
	 332.71 463.95 l
cp p3
np
  335.87 460.68 m
	 338.73 453.77 l
	 338.42 451.55 l
	 335.58 457.71 l
cp p3
np
  338.73 453.77 m
	 341.56 447.24 l
	 341.21 445.61 l
	 338.42 451.55 l
cp p3
np
  341.56 447.24 m
	 344.35 441.12 l
	 343.97 439.98 l
	 341.21 445.61 l
cp p3
np
  344.35 441.12 m
	 347.11 435.43 l
	 346.71 434.70 l
	 343.97 439.98 l
cp p3
np
  347.11 435.43 m
	 349.85 430.19 l
	 349.42 429.79 l
	 346.71 434.70 l
cp p3
np
  349.85 430.19 m
	 352.56 425.40 l
	 352.11 425.28 l
	 349.42 429.79 l
cp p3
np
  352.56 425.40 m
	 355.27 421.05 l
	 354.79 421.17 l
	 352.11 425.28 l
cp p3
np
  277.82 413.64 m
	 280.51 417.13 l
	 281.02 417.46 l
	 278.36 414.15 l
cp p3
np
  280.51 417.13 m
	 283.21 421.05 l
	 283.69 421.17 l
	 281.02 417.46 l
cp p3
np
  283.21 421.05 m
	 285.91 425.40 l
	 286.37 425.28 l
	 283.69 421.17 l
cp p3
np
  285.91 425.40 m
	 288.63 430.19 l
	 289.06 429.79 l
	 286.37 425.28 l
cp p3
np
  288.63 430.19 m
	 291.37 435.43 l
	 291.77 434.70 l
	 289.06 429.79 l
cp p3
np
  291.37 435.43 m
	 294.13 441.12 l
	 294.50 439.98 l
	 291.77 434.70 l
cp p3
np
  294.13 441.12 m
	 296.92 447.24 l
	 297.27 445.61 l
	 294.50 439.98 l
cp p3
np
  296.92 447.24 m
	 299.74 453.77 l
	 300.06 451.55 l
	 297.27 445.61 l
cp p3
np
  264.28 402.94 m
	 267.02 404.24 l
	 267.66 405.27 l
	 264.95 404.04 l
cp p3
np
  267.02 404.24 m
	 269.74 405.87 l
	 270.35 406.81 l
	 267.66 405.27 l
cp p3
np
  269.74 405.87 m
	 272.44 407.95 l
	 273.03 408.76 l
	 270.35 406.81 l
cp p3
np
  272.44 407.95 m
	 275.14 410.58 l
	 275.70 411.24 l
	 273.03 408.76 l
cp p3
np
  275.14 410.58 m
	 277.82 413.64 l
	 278.36 414.15 l
	 275.70 411.24 l
cp p3
np
  299.74 453.77 m
	 302.61 460.68 l
	 302.89 457.71 l
	 300.06 451.55 l
cp p3
np
  302.61 460.68 m
	 305.52 467.86 l
	 305.76 463.95 l
	 302.89 457.71 l
cp p3
np
  305.52 467.86 m
	 308.48 475.13 l
	 308.68 470.04 l
	 305.76 463.95 l
cp p3
np
  361.19 412.92 m
	 363.91 409.74 l
	 363.34 410.58 l
	 360.65 413.64 l
cp p3
np
  353.02 425.16 m
	 355.75 420.62 l
	 355.27 421.05 l
	 352.56 425.40 l
cp p3
np
  355.75 420.62 m
	 358.47 416.54 l
	 357.96 417.13 l
	 355.27 421.05 l
cp p3
np
  358.47 416.54 m
	 361.19 412.92 l
	 360.65 413.64 l
	 357.96 417.13 l
cp p3
np
  372.11 403.11 m
	 374.87 401.75 l
	 374.19 402.94 l
	 371.46 404.24 l
cp p3
np
  363.91 409.74 m
	 366.63 406.99 l
	 366.03 407.95 l
	 363.34 410.58 l
cp p3
np
  366.63 406.99 m
	 369.36 404.81 l
	 368.74 405.87 l
	 366.03 407.95 l
cp p3
np
  369.36 404.81 m
	 372.11 403.11 l
	 371.46 404.24 l
	 368.74 405.87 l
cp p3
np
  302.34 462.75 m
	 305.28 470.77 l
	 305.52 467.86 l
	 302.61 460.68 l
cp p3
np
  305.28 470.77 m
	 308.27 479.19 l
	 308.48 475.13 l
	 305.52 467.86 l
cp p3
np
  308.27 479.19 m
	 311.33 487.78 l
	 311.49 482.12 l
	 308.48 475.13 l
cp p3
np
  311.33 487.78 m
	 314.45 495.92 l
	 314.56 488.07 l
	 311.49 482.12 l
cp p3
np
  314.45 495.92 m
	 317.63 501.73 l
	 317.67 491.72 l
	 314.56 488.07 l
cp p3
np
  317.63 501.73 m
	 320.84 501.73 l
	 320.80 491.72 l
	 317.67 491.72 l
cp p3
np
  320.84 501.73 m
	 324.03 495.92 l
	 323.92 488.07 l
	 320.80 491.72 l
cp p3
np
  324.03 495.92 m
	 327.15 487.78 l
	 326.99 482.12 l
	 323.92 488.07 l
cp p3
np
  327.15 487.78 m
	 330.20 479.19 l
	 330.00 475.13 l
	 326.99 482.12 l
cp p3
np
  330.20 479.19 m
	 333.20 470.77 l
	 332.96 467.86 l
	 330.00 475.13 l
cp p3
np
  333.20 470.77 m
	 336.14 462.75 l
	 335.87 460.68 l
	 332.96 467.86 l
cp p3
np
  336.14 462.75 m
	 339.04 455.22 l
	 338.73 453.77 l
	 335.87 460.68 l
cp p3
np
  339.04 455.22 m
	 341.89 448.19 l
	 341.56 447.24 l
	 338.73 453.77 l
cp p3
np
  341.89 448.19 m
	 344.71 441.68 l
	 344.35 441.12 l
	 341.56 447.24 l
cp p3
np
  344.71 441.68 m
	 347.50 435.68 l
	 347.11 435.43 l
	 344.35 441.12 l
cp p3
np
  347.50 435.68 m
	 350.27 430.17 l
	 349.85 430.19 l
	 347.11 435.43 l
cp p3
np
  350.27 430.17 m
	 353.02 425.16 l
	 352.56 425.40 l
	 349.85 430.19 l
cp p3
np
  274.57 409.74 m
	 277.28 412.92 l
	 277.82 413.64 l
	 275.14 410.58 l
cp p3
np
  277.28 412.92 m
	 280.00 416.54 l
	 280.51 417.13 l
	 277.82 413.64 l
cp p3
np
  280.00 416.54 m
	 282.72 420.62 l
	 283.21 421.05 l
	 280.51 417.13 l
cp p3
np
  282.72 420.62 m
	 285.46 425.16 l
	 285.91 425.40 l
	 283.21 421.05 l
cp p3
np
  285.46 425.16 m
	 288.20 430.17 l
	 288.63 430.19 l
	 285.91 425.40 l
cp p3
np
  288.20 430.17 m
	 290.97 435.68 l
	 291.37 435.43 l
	 288.63 430.19 l
cp p3
np
  290.97 435.68 m
	 293.76 441.68 l
	 294.13 441.12 l
	 291.37 435.43 l
cp p3
np
  293.76 441.68 m
	 296.58 448.19 l
	 296.92 447.24 l
	 294.13 441.12 l
cp p3
np
  296.58 448.19 m
	 299.44 455.22 l
	 299.74 453.77 l
	 296.92 447.24 l
cp p3
np
  263.60 401.75 m
	 266.36 403.11 l
	 267.02 404.24 l
	 264.28 402.94 l
cp p3
np
  266.36 403.11 m
	 269.11 404.81 l
	 269.74 405.87 l
	 267.02 404.24 l
cp p3
np
  269.11 404.81 m
	 271.85 406.99 l
	 272.44 407.95 l
	 269.74 405.87 l
cp p3
np
  271.85 406.99 m
	 274.57 409.74 l
	 275.14 410.58 l
	 272.44 407.95 l
cp p3
np
  299.44 455.22 m
	 302.34 462.75 l
	 302.61 460.68 l
	 299.74 453.77 l
cp p3
np
  350.69 429.66 m
	 353.47 424.50 l
	 353.02 425.16 l
	 350.27 430.17 l
cp p3
np
  356.23 419.84 m
	 358.99 415.66 l
	 358.47 416.54 l
	 355.75 420.62 l
cp p3
np
  358.99 415.66 m
	 361.73 411.94 l
	 361.19 412.92 l
	 358.47 416.54 l
cp p3
np
  361.73 411.94 m
	 364.48 408.68 l
	 363.91 409.74 l
	 361.19 412.92 l
cp p3
np
  353.47 424.50 m
	 356.23 419.84 l
	 355.75 420.62 l
	 353.02 425.16 l
cp p3
np
  367.23 405.86 m
	 369.99 403.62 l
	 369.36 404.81 l
	 366.63 406.99 l
cp p3
np
  369.99 403.62 m
	 372.77 401.87 l
	 372.11 403.11 l
	 369.36 404.81 l
cp p3
np
  372.77 401.87 m
	 375.57 400.48 l
	 374.87 401.75 l
	 372.11 403.11 l
cp p3
np
  364.48 408.68 m
	 367.23 405.86 l
	 366.63 406.99 l
	 363.91 409.74 l
cp p3
np
  299.15 455.65 m
	 302.08 463.59 l
	 302.34 462.75 l
	 299.44 455.22 l
cp p3
np
  302.08 463.59 m
	 305.06 472.16 l
	 305.28 470.77 l
	 302.34 462.75 l
cp p3
np
  305.06 472.16 m
	 308.09 481.37 l
	 308.27 479.19 l
	 305.28 470.77 l
cp p3
np
  308.09 481.37 m
	 311.19 491.23 l
	 311.33 487.78 l
	 308.27 479.19 l
cp p3
np
  311.19 491.23 m
	 314.35 501.62 l
	 314.45 495.92 l
	 311.33 487.78 l
cp p3
np
  314.35 501.62 m
	 317.59 511.65 l
	 317.63 501.73 l
	 314.45 495.92 l
cp p3
np
  317.59 511.65 m
	 320.89 511.65 l
	 320.84 501.73 l
	 317.63 501.73 l
cp p3
np
  320.89 511.65 m
	 324.13 501.62 l
	 324.03 495.92 l
	 320.84 501.73 l
cp p3
np
  324.13 501.62 m
	 327.29 491.23 l
	 327.15 487.78 l
	 324.03 495.92 l
cp p3
np
  327.29 491.23 m
	 330.38 481.37 l
	 330.20 479.19 l
	 327.15 487.78 l
cp p3
np
  330.38 481.37 m
	 333.42 472.16 l
	 333.20 470.77 l
	 330.20 479.19 l
cp p3
np
  333.42 472.16 m
	 336.40 463.59 l
	 336.14 462.75 l
	 333.20 470.77 l
cp p3
np
  336.40 463.59 m
	 339.33 455.65 l
	 339.04 455.22 l
	 336.14 462.75 l
cp p3
np
  339.33 455.65 m
	 342.22 448.31 l
	 341.89 448.19 l
	 339.04 455.22 l
cp p3
np
  342.22 448.31 m
	 345.07 441.55 l
	 344.71 441.68 l
	 341.89 448.19 l
cp p3
np
  345.07 441.55 m
	 347.89 435.34 l
	 347.50 435.68 l
	 344.71 441.68 l
cp p3
np
  347.89 435.34 m
	 350.69 429.66 l
	 350.27 430.17 l
	 347.50 435.68 l
cp p3
np
  265.70 401.87 m
	 268.48 403.62 l
	 269.11 404.81 l
	 266.36 403.11 l
cp p3
np
  268.48 403.62 m
	 271.25 405.86 l
	 271.85 406.99 l
	 269.11 404.81 l
cp p3
np
  271.25 405.86 m
	 274.00 408.68 l
	 274.57 409.74 l
	 271.85 406.99 l
cp p3
np
  274.00 408.68 m
	 276.74 411.94 l
	 277.28 412.92 l
	 274.57 409.74 l
cp p3
np
  276.74 411.94 m
	 279.49 415.66 l
	 280.00 416.54 l
	 277.28 412.92 l
cp p3
np
  279.49 415.66 m
	 282.24 419.84 l
	 282.72 420.62 l
	 280.00 416.54 l
cp p3
np
  282.24 419.84 m
	 285.01 424.50 l
	 285.46 425.16 l
	 282.72 420.62 l
cp p3
np
  285.01 424.50 m
	 287.79 429.66 l
	 288.20 430.17 l
	 285.46 425.16 l
cp p3
np
  287.79 429.66 m
	 290.58 435.34 l
	 290.97 435.68 l
	 288.20 430.17 l
cp p3
np
  290.58 435.34 m
	 293.41 441.55 l
	 293.76 441.68 l
	 290.97 435.68 l
cp p3
np
  293.41 441.55 m
	 296.26 448.31 l
	 296.58 448.19 l
	 293.76 441.68 l
cp p3
np
  296.26 448.31 m
	 299.15 455.65 l
	 299.44 455.22 l
	 296.58 448.19 l
cp p3
np
  262.91 400.48 m
	 265.70 401.87 l
	 266.36 403.11 l
	 263.60 401.75 l
cp p3
np
  342.52 447.50 m
	 345.41 440.65 l
	 345.07 441.55 l
	 342.22 448.31 l
cp p3
np
  345.41 440.65 m
	 348.27 434.37 l
	 347.89 435.34 l
	 345.07 441.55 l
cp p3
np
  348.27 434.37 m
	 351.10 428.63 l
	 350.69 429.66 l
	 347.89 435.34 l
cp p3
np
  351.10 428.63 m
	 353.91 423.40 l
	 353.47 424.50 l
	 350.69 429.66 l
cp p3
np
  353.91 423.40 m
	 356.71 418.69 l
	 356.23 419.84 l
	 353.47 424.50 l
cp p3
np
  356.71 418.69 m
	 359.49 414.46 l
	 358.99 415.66 l
	 356.23 419.84 l
cp p3
np
  359.49 414.46 m
	 362.27 410.70 l
	 361.73 411.94 l
	 358.99 415.66 l
cp p3
np
  362.27 410.70 m
	 365.05 407.40 l
	 364.48 408.68 l
	 361.73 411.94 l
cp p3
np
  365.05 407.40 m
	 367.83 404.55 l
	 367.23 405.86 l
	 364.48 408.68 l
cp p3
np
  367.83 404.55 m
	 370.63 402.29 l
	 369.99 403.62 l
	 367.23 405.86 l
cp p3
np
  370.63 402.29 m
	 373.45 400.52 l
	 372.77 401.87 l
	 369.99 403.62 l
cp p3
np
  373.45 400.52 m
	 376.28 399.11 l
	 375.57 400.48 l
	 372.77 401.87 l
cp p3
np
  295.95 447.50 m
	 298.88 454.93 l
	 299.15 455.65 l
	 296.26 448.31 l
cp p3
np
  298.88 454.93 m
	 301.85 462.97 l
	 302.08 463.59 l
	 299.15 455.65 l
cp p3
np
  301.85 462.97 m
	 304.86 471.65 l
	 305.06 472.16 l
	 302.08 463.59 l
cp p3
np
  304.86 471.65 m
	 307.94 480.99 l
	 308.09 481.37 l
	 305.06 472.16 l
cp p3
np
  307.94 480.99 m
	 311.07 490.97 l
	 311.19 491.23 l
	 308.09 481.37 l
cp p3
np
  311.07 490.97 m
	 314.28 501.51 l
	 314.35 501.62 l
	 311.19 491.23 l
cp p3
np
  314.28 501.51 m
	 317.57 511.68 l
	 317.59 511.65 l
	 314.35 501.62 l
cp p3
np
  317.57 511.68 m
	 320.91 511.68 l
	 320.89 511.65 l
	 317.59 511.65 l
cp p3
np
  320.91 511.68 m
	 324.20 501.51 l
	 324.13 501.62 l
	 320.89 511.65 l
cp p3
np
  324.20 501.51 m
	 327.40 490.97 l
	 327.29 491.23 l
	 324.13 501.62 l
cp p3
np
  327.40 490.97 m
	 330.54 480.99 l
	 330.38 481.37 l
	 327.29 491.23 l
cp p3
np
  330.54 480.99 m
	 333.61 471.65 l
	 333.42 472.16 l
	 330.38 481.37 l
cp p3
np
  333.61 471.65 m
	 336.63 462.97 l
	 336.40 463.59 l
	 333.42 472.16 l
cp p3
np
  336.63 462.97 m
	 339.60 454.93 l
	 339.33 455.65 l
	 336.40 463.59 l
cp p3
np
  339.60 454.93 m
	 342.52 447.50 l
	 342.22 448.31 l
	 339.33 455.65 l
cp p3
np
  262.20 399.11 m
	 265.03 400.52 l
	 265.70 401.87 l
	 262.91 400.48 l
cp p3
np
  265.03 400.52 m
	 267.84 402.29 l
	 268.48 403.62 l
	 265.70 401.87 l
cp p3
np
  267.84 402.29 m
	 270.64 404.55 l
	 271.25 405.86 l
	 268.48 403.62 l
cp p3
np
  270.64 404.55 m
	 273.42 407.40 l
	 274.00 408.68 l
	 271.25 405.86 l
cp p3
np
  273.42 407.40 m
	 276.20 410.70 l
	 276.74 411.94 l
	 274.00 408.68 l
cp p3
np
  276.20 410.70 m
	 278.98 414.46 l
	 279.49 415.66 l
	 276.74 411.94 l
cp p3
np
  278.98 414.46 m
	 281.77 418.69 l
	 282.24 419.84 l
	 279.49 415.66 l
cp p3
np
  281.77 418.69 m
	 284.56 423.40 l
	 285.01 424.50 l
	 282.24 419.84 l
cp p3
np
  284.56 423.40 m
	 287.38 428.63 l
	 287.79 429.66 l
	 285.01 424.50 l
cp p3
np
  287.38 428.63 m
	 290.21 434.37 l
	 290.58 435.34 l
	 287.79 429.66 l
cp p3
np
  290.21 434.37 m
	 293.07 440.65 l
	 293.41 441.55 l
	 290.58 435.34 l
cp p3
np
  293.07 440.65 m
	 295.95 447.50 l
	 296.26 448.31 l
	 293.41 441.55 l
cp p3
np
  374.13 399.04 m
	 377.00 397.64 l
	 376.28 399.11 l
	 373.45 400.52 l
cp p3
np
  339.85 453.00 m
	 342.81 445.71 l
	 342.52 447.50 l
	 339.60 454.93 l
cp p3
np
  342.81 445.71 m
	 345.74 438.96 l
	 345.41 440.65 l
	 342.52 447.50 l
cp p3
np
  345.74 438.96 m
	 348.63 432.74 l
	 348.27 434.37 l
	 345.41 440.65 l
cp p3
np
  348.63 432.74 m
	 351.50 427.03 l
	 351.10 428.63 l
	 348.27 434.37 l
cp p3
np
  351.50 427.03 m
	 354.35 421.84 l
	 353.91 423.40 l
	 351.10 428.63 l
cp p3
np
  354.35 421.84 m
	 357.18 417.14 l
	 356.71 418.69 l
	 353.91 423.40 l
cp p3
np
  357.18 417.14 m
	 360.00 412.93 l
	 359.49 414.46 l
	 356.71 418.69 l
cp p3
np
  360.00 412.93 m
	 362.82 409.18 l
	 362.27 410.70 l
	 359.49 414.46 l
cp p3
np
  362.82 409.18 m
	 365.63 405.89 l
	 365.05 407.40 l
	 362.27 410.70 l
cp p3
np
  365.63 405.89 m
	 368.45 403.05 l
	 367.83 404.55 l
	 365.05 407.40 l
cp p3
np
  368.45 403.05 m
	 371.28 400.81 l
	 370.63 402.29 l
	 367.83 404.55 l
cp p3
np
  371.28 400.81 m
	 374.13 399.04 l
	 373.45 400.52 l
	 370.63 402.29 l
cp p3
np
  286.97 427.03 m
	 289.84 432.74 l
	 290.21 434.37 l
	 287.38 428.63 l
cp p3
np
  289.84 432.74 m
	 292.74 438.96 l
	 293.07 440.65 l
	 290.21 434.37 l
cp p3
np
  292.74 438.96 m
	 295.67 445.71 l
	 295.95 447.50 l
	 293.07 440.65 l
cp p3
np
  295.67 445.71 m
	 298.63 453.00 l
	 298.88 454.93 l
	 295.95 447.50 l
cp p3
np
  298.63 453.00 m
	 301.64 460.83 l
	 301.85 462.97 l
	 298.88 454.93 l
cp p3
np
  301.64 460.83 m
	 304.70 469.16 l
	 304.86 471.65 l
	 301.85 462.97 l
cp p3
np
  304.70 469.16 m
	 307.81 477.92 l
	 307.94 480.99 l
	 304.86 471.65 l
cp p3
np
  307.81 477.92 m
	 310.99 486.87 l
	 311.07 490.97 l
	 307.94 480.99 l
cp p3
np
  310.99 486.87 m
	 314.24 495.34 l
	 314.28 501.51 l
	 311.07 490.97 l
cp p3
np
  314.24 495.34 m
	 317.56 501.40 l
	 317.57 511.68 l
	 314.28 501.51 l
cp p3
np
  317.56 501.40 m
	 320.91 501.40 l
	 320.91 511.68 l
	 317.57 511.68 l
cp p3
np
  320.91 501.40 m
	 324.23 495.34 l
	 324.20 501.51 l
	 320.91 511.68 l
cp p3
np
  324.23 495.34 m
	 327.48 486.87 l
	 327.40 490.97 l
	 324.20 501.51 l
cp p3
np
  327.48 486.87 m
	 330.66 477.92 l
	 330.54 480.99 l
	 327.40 490.97 l
cp p3
np
  330.66 477.92 m
	 333.78 469.16 l
	 333.61 471.65 l
	 330.54 480.99 l
cp p3
np
  333.78 469.16 m
	 336.84 460.83 l
	 336.63 462.97 l
	 333.61 471.65 l
cp p3
np
  336.84 460.83 m
	 339.85 453.00 l
	 339.60 454.93 l
	 336.63 462.97 l
cp p3
np
  270.03 403.05 m
	 272.84 405.89 l
	 273.42 407.40 l
	 270.64 404.55 l
cp p3
np
  261.48 397.64 m
	 264.34 399.04 l
	 265.03 400.52 l
	 262.20 399.11 l
cp p3
np
  264.34 399.04 m
	 267.19 400.81 l
	 267.84 402.29 l
	 265.03 400.52 l
cp p3
np
  267.19 400.81 m
	 270.03 403.05 l
	 270.64 404.55 l
	 267.84 402.29 l
cp p3
np
  281.29 417.14 m
	 284.13 421.84 l
	 284.56 423.40 l
	 281.77 418.69 l
cp p3
np
  272.84 405.89 m
	 275.66 409.18 l
	 276.20 410.70 l
	 273.42 407.40 l
cp p3
np
  275.66 409.18 m
	 278.47 412.93 l
	 278.98 414.46 l
	 276.20 410.70 l
cp p3
np
  278.47 412.93 m
	 281.29 417.14 l
	 281.77 418.69 l
	 278.98 414.46 l
cp p3
np
  284.13 421.84 m
	 286.97 427.03 l
	 287.38 428.63 l
	 284.56 423.40 l
cp p3
np
  337.02 457.30 m
	 340.07 449.95 l
	 339.85 453.00 l
	 336.84 460.83 l
cp p3
np
  366.21 404.15 m
	 369.07 401.37 l
	 368.45 403.05 l
	 365.63 405.89 l
cp p3
np
  369.07 401.37 m
	 371.94 399.17 l
	 371.28 400.81 l
	 368.45 403.05 l
cp p3
np
  371.94 399.17 m
	 374.83 397.45 l
	 374.13 399.04 l
	 371.28 400.81 l
cp p3
np
  374.83 397.45 m
	 377.73 396.08 l
	 377.00 397.64 l
	 374.13 399.04 l
cp p3
np
  340.07 449.95 m
	 343.08 442.99 l
	 342.81 445.71 l
	 339.85 453.00 l
cp p3
np
  343.08 442.99 m
	 346.05 436.49 l
	 345.74 438.96 l
	 342.81 445.71 l
cp p3
np
  346.05 436.49 m
	 348.98 430.46 l
	 348.63 432.74 l
	 345.74 438.96 l
cp p3
np
  348.98 430.46 m
	 351.89 424.90 l
	 351.50 427.03 l
	 348.63 432.74 l
cp p3
np
  351.89 424.90 m
	 354.78 419.82 l
	 354.35 421.84 l
	 351.50 427.03 l
cp p3
np
  354.78 419.82 m
	 357.65 415.21 l
	 357.18 417.14 l
	 354.35 421.84 l
cp p3
np
  357.65 415.21 m
	 360.51 411.07 l
	 360.00 412.93 l
	 357.18 417.14 l
cp p3
np
  360.51 411.07 m
	 363.36 407.38 l
	 362.82 409.18 l
	 360.00 412.93 l
cp p3
np
  363.36 407.38 m
	 366.21 404.15 l
	 365.63 405.89 l
	 362.82 409.18 l
cp p3
np
  283.70 419.82 m
	 286.58 424.90 l
	 286.97 427.03 l
	 284.13 421.84 l
cp p3
np
  286.58 424.90 m
	 289.49 430.46 l
	 289.84 432.74 l
	 286.97 427.03 l
cp p3
np
  289.49 430.46 m
	 292.43 436.49 l
	 292.74 438.96 l
	 289.84 432.74 l
cp p3
np
  292.43 436.49 m
	 295.40 442.99 l
	 295.67 445.71 l
	 292.74 438.96 l
cp p3
np
  295.40 442.99 m
	 298.40 449.95 l
	 298.63 453.00 l
	 295.67 445.71 l
cp p3
np
  298.40 449.95 m
	 301.45 457.30 l
	 301.64 460.83 l
	 298.63 453.00 l
cp p3
np
  301.45 457.30 m
	 304.56 464.95 l
	 304.70 469.16 l
	 301.64 460.83 l
cp p3
np
  304.56 464.95 m
	 307.71 472.71 l
	 307.81 477.92 l
	 304.70 469.16 l
cp p3
np
  307.71 472.71 m
	 310.94 480.17 l
	 310.99 486.87 l
	 307.81 477.92 l
cp p3
np
  310.94 480.17 m
	 314.22 486.54 l
	 314.24 495.34 l
	 310.99 486.87 l
cp p3
np
  314.22 486.54 m
	 317.56 490.44 l
	 317.56 501.40 l
	 314.24 495.34 l
cp p3
np
  317.56 490.44 m
	 320.92 490.44 l
	 320.91 501.40 l
	 317.56 501.40 l
cp p3
np
  320.92 490.44 m
	 324.26 486.54 l
	 324.23 495.34 l
	 320.91 501.40 l
cp p3
np
  324.26 486.54 m
	 327.54 480.17 l
	 327.48 486.87 l
	 324.23 495.34 l
cp p3
np
  327.54 480.17 m
	 330.76 472.71 l
	 330.66 477.92 l
	 327.48 486.87 l
cp p3
np
  330.76 472.71 m
	 333.92 464.95 l
	 333.78 469.16 l
	 330.66 477.92 l
cp p3
np
  333.92 464.95 m
	 337.02 457.30 l
	 336.84 460.83 l
	 333.78 469.16 l
cp p3
np
  263.64 397.45 m
	 266.53 399.17 l
	 267.19 400.81 l
	 264.34 399.04 l
cp p3
np
  266.53 399.17 m
	 269.41 401.37 l
	 270.03 403.05 l
	 267.19 400.81 l
cp p3
np
  269.41 401.37 m
	 272.26 404.15 l
	 272.84 405.89 l
	 270.03 403.05 l
cp p3
np
  260.74 396.08 m
	 263.64 397.45 l
	 264.34 399.04 l
	 261.48 397.64 l
cp p3
np
  275.11 407.38 m
	 277.97 411.07 l
	 278.47 412.93 l
	 275.66 409.18 l
cp p3
np
  277.97 411.07 m
	 280.83 415.21 l
	 281.29 417.14 l
	 278.47 412.93 l
cp p3
np
  280.83 415.21 m
	 283.70 419.82 l
	 284.13 421.84 l
	 281.29 417.14 l
cp p3
np
  272.26 404.15 m
	 275.11 407.38 l
	 275.66 409.18 l
	 272.84 405.89 l
cp p3
np
  330.84 466.12 m
	 334.04 459.46 l
	 333.92 464.95 l
	 330.76 472.71 l
cp p3
np
  334.04 459.46 m
	 337.19 452.64 l
	 337.02 457.30 l
	 333.92 464.95 l
cp p3
np
  337.19 452.64 m
	 340.28 445.92 l
	 340.07 449.95 l
	 337.02 457.30 l
cp p3
np
  363.91 405.32 m
	 366.80 402.18 l
	 366.21 404.15 l
	 363.36 407.38 l
cp p3
np
  366.80 402.18 m
	 369.69 399.50 l
	 369.07 401.37 l
	 366.21 404.15 l
cp p3
np
  369.69 399.50 m
	 372.61 397.40 l
	 371.94 399.17 l
	 369.07 401.37 l
cp p3
np
  372.61 397.40 m
	 375.54 395.74 l
	 374.83 397.45 l
	 371.94 399.17 l
cp p3
np
  375.54 395.74 m
	 378.48 394.41 l
	 377.73 396.08 l
	 374.83 397.45 l
cp p3
np
  340.28 445.92 m
	 343.33 439.45 l
	 343.08 442.99 l
	 340.07 449.95 l
cp p3
np
  343.33 439.45 m
	 346.34 433.32 l
	 346.05 436.49 l
	 343.08 442.99 l
cp p3
np
  346.34 433.32 m
	 349.32 427.58 l
	 348.98 430.46 l
	 346.05 436.49 l
cp p3
np
  349.32 427.58 m
	 352.27 422.26 l
	 351.89 424.90 l
	 348.98 430.46 l
cp p3
np
  352.27 422.26 m
	 355.20 417.37 l
	 354.78 419.82 l
	 351.89 424.90 l
cp p3
np
  355.20 417.37 m
	 358.11 412.91 l
	 357.65 415.21 l
	 354.78 419.82 l
cp p3
np
  358.11 412.91 m
	 361.01 408.90 l
	 360.51 411.07 l
	 357.65 415.21 l
cp p3
np
  361.01 408.90 m
	 363.91 405.32 l
	 363.36 407.38 l
	 360.51 411.07 l
cp p3
np
  280.36 412.91 m
	 283.27 417.37 l
	 283.70 419.82 l
	 280.83 415.21 l
cp p3
np
  283.27 417.37 m
	 286.20 422.26 l
	 286.58 424.90 l
	 283.70 419.82 l
cp p3
np
  286.20 422.26 m
	 289.15 427.58 l
	 289.49 430.46 l
	 286.58 424.90 l
cp p3
np
  289.15 427.58 m
	 292.13 433.32 l
	 292.43 436.49 l
	 289.49 430.46 l
cp p3
np
  292.13 433.32 m
	 295.14 439.45 l
	 295.40 442.99 l
	 292.43 436.49 l
cp p3
np
  295.14 439.45 m
	 298.19 445.92 l
	 298.40 449.95 l
	 295.40 442.99 l
cp p3
np
  298.19 445.92 m
	 301.29 452.64 l
	 301.45 457.30 l
	 298.40 449.95 l
cp p3
np
  301.29 452.64 m
	 304.43 459.46 l
	 304.56 464.95 l
	 301.45 457.30 l
cp p3
np
  304.43 459.46 m
	 307.63 466.12 l
	 307.71 472.71 l
	 304.56 464.95 l
cp p3
np
  307.63 466.12 m
	 310.89 472.19 l
	 310.94 480.17 l
	 307.71 472.71 l
cp p3
np
  310.89 472.19 m
	 314.20 477.01 l
	 314.22 486.54 l
	 310.94 480.17 l
cp p3
np
  314.20 477.01 m
	 317.55 479.75 l
	 317.56 490.44 l
	 314.22 486.54 l
cp p3
np
  317.55 479.75 m
	 320.92 479.75 l
	 320.92 490.44 l
	 317.56 490.44 l
cp p3
np
  320.92 479.75 m
	 324.28 477.01 l
	 324.26 486.54 l
	 320.92 490.44 l
cp p3
np
  324.28 477.01 m
	 327.59 472.19 l
	 327.54 480.17 l
	 324.26 486.54 l
cp p3
np
  327.59 472.19 m
	 330.84 466.12 l
	 330.76 472.71 l
	 327.54 480.17 l
cp p3
np
  259.99 394.41 m
	 262.93 395.74 l
	 263.64 397.45 l
	 260.74 396.08 l
cp p3
np
  262.93 395.74 m
	 265.87 397.40 l
	 266.53 399.17 l
	 263.64 397.45 l
cp p3
np
  265.87 397.40 m
	 268.78 399.50 l
	 269.41 401.37 l
	 266.53 399.17 l
cp p3
np
  268.78 399.50 m
	 271.68 402.18 l
	 272.26 404.15 l
	 269.41 401.37 l
cp p3
np
  271.68 402.18 m
	 274.57 405.32 l
	 275.11 407.38 l
	 272.26 404.15 l
cp p3
np
  274.57 405.32 m
	 277.46 408.90 l
	 277.97 411.07 l
	 275.11 407.38 l
cp p3
np
  277.46 408.90 m
	 280.36 412.91 l
	 280.83 415.21 l
	 277.97 411.07 l
cp p3
np
  337.34 447.15 m
	 340.48 441.13 l
	 340.28 445.92 l
	 337.19 452.64 l
cp p3
np
  327.63 463.67 m
	 330.92 458.74 l
	 330.84 466.12 l
	 327.59 472.19 l
cp p3
np
  330.92 458.74 m
	 334.16 453.11 l
	 334.04 459.46 l
	 330.84 466.12 l
cp p3
np
  334.16 453.11 m
	 337.34 447.15 l
	 337.19 452.64 l
	 334.04 459.46 l
cp p3
np
  361.52 406.44 m
	 364.45 403.02 l
	 363.91 405.32 l
	 361.01 408.90 l
cp p3
np
  364.45 403.02 m
	 367.39 400.01 l
	 366.80 402.18 l
	 363.91 405.32 l
cp p3
np
  367.39 400.01 m
	 370.33 397.48 l
	 369.69 399.50 l
	 366.80 402.18 l
cp p3
np
  370.33 397.48 m
	 373.29 395.50 l
	 372.61 397.40 l
	 369.69 399.50 l
cp p3
np
  373.29 395.50 m
	 376.26 393.92 l
	 375.54 395.74 l
	 372.61 397.40 l
cp p3
np
  376.26 393.92 m
	 379.25 392.65 l
	 378.48 394.41 l
	 375.54 395.74 l
cp p3
np
  340.48 441.13 m
	 343.58 435.23 l
	 343.33 439.45 l
	 340.28 445.92 l
cp p3
np
  343.58 435.23 m
	 346.63 429.55 l
	 346.34 433.32 l
	 343.33 439.45 l
cp p3
np
  346.63 429.55 m
	 349.65 424.18 l
	 349.32 427.58 l
	 346.34 433.32 l
cp p3
np
  349.65 424.18 m
	 352.65 419.16 l
	 352.27 422.26 l
	 349.32 427.58 l
cp p3
np
  352.65 419.16 m
	 355.62 414.52 l
	 355.20 417.37 l
	 352.27 422.26 l
cp p3
np
  355.62 414.52 m
	 358.57 410.28 l
	 358.11 412.91 l
	 355.20 417.37 l
cp p3
np
  358.57 410.28 m
	 361.52 406.44 l
	 361.01 408.90 l
	 358.11 412.91 l
cp p3
np
  274.02 403.02 m
	 276.96 406.44 l
	 277.46 408.90 l
	 274.57 405.32 l
cp p3
np
  276.96 406.44 m
	 279.90 410.28 l
	 280.36 412.91 l
	 277.46 408.90 l
cp p3
np
  279.90 410.28 m
	 282.86 414.52 l
	 283.27 417.37 l
	 280.36 412.91 l
cp p3
np
  282.86 414.52 m
	 285.83 419.16 l
	 286.20 422.26 l
	 283.27 417.37 l
cp p3
np
  285.83 419.16 m
	 288.82 424.18 l
	 289.15 427.58 l
	 286.20 422.26 l
cp p3
np
  288.82 424.18 m
	 291.85 429.55 l
	 292.13 433.32 l
	 289.15 427.58 l
cp p3
np
  291.85 429.55 m
	 294.90 435.23 l
	 295.14 439.45 l
	 292.13 433.32 l
cp p3
np
  294.90 435.23 m
	 297.99 441.13 l
	 298.19 445.92 l
	 295.14 439.45 l
cp p3
np
  297.99 441.13 m
	 301.13 447.15 l
	 301.29 452.64 l
	 298.19 445.92 l
cp p3
np
  301.13 447.15 m
	 304.32 453.11 l
	 304.43 459.46 l
	 301.29 452.64 l
cp p3
np
  304.32 453.11 m
	 307.56 458.74 l
	 307.63 466.12 l
	 304.43 459.46 l
cp p3
np
  307.56 458.74 m
	 310.85 463.67 l
	 310.89 472.19 l
	 307.63 466.12 l
cp p3
np
  310.85 463.67 m
	 314.18 467.41 l
	 314.20 477.01 l
	 310.89 472.19 l
cp p3
np
  314.18 467.41 m
	 317.55 469.46 l
	 317.55 479.75 l
	 314.20 477.01 l
cp p3
np
  317.55 469.46 m
	 320.93 469.46 l
	 320.92 479.75 l
	 317.55 479.75 l
cp p3
np
  320.93 469.46 m
	 324.30 467.41 l
	 324.28 477.01 l
	 320.92 479.75 l
cp p3
np
  324.30 467.41 m
	 327.63 463.67 l
	 327.59 472.19 l
	 324.28 477.01 l
cp p3
np
  268.15 397.48 m
	 271.09 400.01 l
	 271.68 402.18 l
	 268.78 399.50 l
cp p3
np
  259.23 392.65 m
	 262.21 393.92 l
	 262.93 395.74 l
	 259.99 394.41 l
cp p3
np
  262.21 393.92 m
	 265.19 395.50 l
	 265.87 397.40 l
	 262.93 395.74 l
cp p3
np
  265.19 395.50 m
	 268.15 397.48 l
	 268.78 399.50 l
	 265.87 397.40 l
cp p3
np
  271.09 400.01 m
	 274.02 403.02 l
	 274.57 405.32 l
	 271.68 402.18 l
cp p3
np
  324.32 458.00 m
	 327.67 455.03 l
	 327.63 463.67 l
	 324.30 467.41 l
cp p3
np
  330.99 451.00 m
	 334.26 446.26 l
	 334.16 453.11 l
	 330.92 458.74 l
cp p3
np
  334.26 446.26 m
	 337.49 441.10 l
	 337.34 447.15 l
	 334.16 453.11 l
cp p3
np
  337.49 441.10 m
	 340.67 435.78 l
	 340.48 441.13 l
	 337.34 447.15 l
cp p3
np
  327.67 455.03 m
	 330.99 451.00 l
	 330.92 458.74 l
	 327.63 463.67 l
cp p3
np
  356.03 411.33 m
	 359.03 407.34 l
	 358.57 410.28 l
	 355.62 414.52 l
cp p3
np
  359.03 407.34 m
	 362.02 403.72 l
	 361.52 406.44 l
	 358.57 410.28 l
cp p3
np
  362.02 403.72 m
	 365.00 400.49 l
	 364.45 403.02 l
	 361.52 406.44 l
cp p3
np
  365.00 400.49 m
	 367.98 397.64 l
	 367.39 400.01 l
	 364.45 403.02 l
cp p3
np
  367.98 397.64 m
	 370.98 395.32 l
	 370.33 397.48 l
	 367.39 400.01 l
cp p3
np
  370.98 395.32 m
	 373.98 393.48 l
	 373.29 395.50 l
	 370.33 397.48 l
cp p3
np
  373.98 393.48 m
	 377.00 392.00 l
	 376.26 393.92 l
	 373.29 395.50 l
cp p3
np
  377.00 392.00 m
	 380.03 390.80 l
	 379.25 392.65 l
	 376.26 393.92 l
cp p3
np
  340.67 435.78 m
	 343.81 430.47 l
	 343.58 435.23 l
	 340.48 441.13 l
cp p3
np
  343.81 430.47 m
	 346.91 425.29 l
	 346.63 429.55 l
	 343.58 435.23 l
cp p3
np
  346.91 425.29 m
	 349.98 420.34 l
	 349.65 424.18 l
	 346.63 429.55 l
cp p3
np
  349.98 420.34 m
	 353.02 415.67 l
	 352.65 419.16 l
	 349.65 424.18 l
cp p3
np
  353.02 415.67 m
	 356.03 411.33 l
	 355.62 414.52 l
	 352.65 419.16 l
cp p3
np
  270.49 397.64 m
	 273.47 400.49 l
	 274.02 403.02 l
	 271.09 400.01 l
cp p3
np
  273.47 400.49 m
	 276.45 403.72 l
	 276.96 406.44 l
	 274.02 403.02 l
cp p3
np
  276.45 403.72 m
	 279.44 407.34 l
	 279.90 410.28 l
	 276.96 406.44 l
cp p3
np
  279.44 407.34 m
	 282.44 411.33 l
	 282.86 414.52 l
	 279.90 410.28 l
cp p3
np
  282.44 411.33 m
	 285.46 415.67 l
	 285.83 419.16 l
	 282.86 414.52 l
cp p3
np
  285.46 415.67 m
	 288.50 420.34 l
	 288.82 424.18 l
	 285.83 419.16 l
cp p3
np
  288.50 420.34 m
	 291.57 425.29 l
	 291.85 429.55 l
	 288.82 424.18 l
cp p3
np
  291.57 425.29 m
	 294.67 430.47 l
	 294.90 435.23 l
	 291.85 429.55 l
cp p3
np
  294.67 430.47 m
	 297.81 435.78 l
	 297.99 441.13 l
	 294.90 435.23 l
cp p3
np
  297.81 435.78 m
	 300.99 441.10 l
	 301.13 447.15 l
	 297.99 441.13 l
cp p3
np
  300.99 441.10 m
	 304.21 446.26 l
	 304.32 453.11 l
	 301.13 447.15 l
cp p3
np
  304.21 446.26 m
	 307.48 451.00 l
	 307.56 458.74 l
	 304.32 453.11 l
cp p3
np
  307.48 451.00 m
	 310.80 455.03 l
	 310.85 463.67 l
	 307.56 458.74 l
cp p3
np
  310.80 455.03 m
	 314.16 458.00 l
	 314.18 467.41 l
	 310.85 463.67 l
cp p3
np
  314.16 458.00 m
	 317.54 459.59 l
	 317.55 469.46 l
	 314.18 467.41 l
cp p3
np
  317.54 459.59 m
	 320.93 459.59 l
	 320.93 469.46 l
	 317.55 469.46 l
cp p3
np
  320.93 459.59 m
	 324.32 458.00 l
	 324.30 467.41 l
	 320.93 469.46 l
cp p3
np
  261.47 392.00 m
	 264.49 393.48 l
	 265.19 395.50 l
	 262.21 393.92 l
cp p3
np
  264.49 393.48 m
	 267.50 395.32 l
	 268.15 397.48 l
	 265.19 395.50 l
cp p3
np
  267.50 395.32 m
	 270.49 397.64 l
	 271.09 400.01 l
	 268.15 397.48 l
cp p3
np
  258.44 390.80 m
	 261.47 392.00 l
	 262.21 393.92 l
	 259.23 392.65 l
cp p3
np
  317.53 450.15 m
	 320.94 450.15 l
	 320.93 459.59 l
	 317.54 459.59 l
cp p3
np
  320.94 450.15 m
	 324.34 448.88 l
	 324.32 458.00 l
	 320.93 459.59 l
cp p3
np
  324.34 448.88 m
	 327.72 446.48 l
	 327.67 455.03 l
	 324.32 458.00 l
cp p3
np
  327.72 446.48 m
	 331.06 443.15 l
	 330.99 451.00 l
	 327.67 455.03 l
cp p3
np
  331.06 443.15 m
	 334.37 439.16 l
	 334.26 446.26 l
	 330.99 451.00 l
cp p3
np
  334.37 439.16 m
	 337.63 434.72 l
	 337.49 441.10 l
	 334.26 446.26 l
cp p3
np
  337.63 434.72 m
	 340.86 430.06 l
	 340.67 435.78 l
	 337.49 441.10 l
cp p3
np
  353.38 411.87 m
	 356.45 407.85 l
	 356.03 411.33 l
	 353.02 415.67 l
cp p3
np
  356.45 407.85 m
	 359.50 404.15 l
	 359.03 407.34 l
	 356.03 411.33 l
cp p3
np
  359.50 404.15 m
	 362.53 400.78 l
	 362.02 403.72 l
	 359.03 407.34 l
cp p3
np
  362.53 400.78 m
	 365.56 397.77 l
	 365.00 400.49 l
	 362.02 403.72 l
cp p3
np
  365.56 397.77 m
	 368.59 395.14 l
	 367.98 397.64 l
	 365.00 400.49 l
cp p3
np
  368.59 395.14 m
	 371.64 393.04 l
	 370.98 395.32 l
	 367.98 397.64 l
cp p3
np
  371.64 393.04 m
	 374.69 391.35 l
	 373.98 393.48 l
	 370.98 395.32 l
cp p3
np
  374.69 391.35 m
	 377.76 389.98 l
	 377.00 392.00 l
	 373.98 393.48 l
cp p3
np
  377.76 389.98 m
	 380.83 388.86 l
	 380.03 390.80 l
	 377.00 392.00 l
cp p3
np
  340.86 430.06 m
	 344.04 425.33 l
	 343.81 430.47 l
	 340.67 435.78 l
cp p3
np
  344.04 425.33 m
	 347.18 420.67 l
	 346.91 425.29 l
	 343.81 430.47 l
cp p3
np
  347.18 420.67 m
	 350.30 416.16 l
	 349.98 420.34 l
	 346.91 425.29 l
cp p3
np
  350.30 416.16 m
	 353.38 411.87 l
	 353.02 415.67 l
	 349.98 420.34 l
cp p3
np
  266.84 393.04 m
	 269.88 395.14 l
	 270.49 397.64 l
	 267.50 395.32 l
cp p3
np
  269.88 395.14 m
	 272.91 397.77 l
	 273.47 400.49 l
	 270.49 397.64 l
cp p3
np
  272.91 397.77 m
	 275.94 400.78 l
	 276.45 403.72 l
	 273.47 400.49 l
cp p3
np
  275.94 400.78 m
	 278.98 404.15 l
	 279.44 407.34 l
	 276.45 403.72 l
cp p3
np
  278.98 404.15 m
	 282.03 407.85 l
	 282.44 411.33 l
	 279.44 407.34 l
cp p3
np
  282.03 407.85 m
	 285.09 411.87 l
	 285.46 415.67 l
	 282.44 411.33 l
cp p3
np
  285.09 411.87 m
	 288.18 416.16 l
	 288.50 420.34 l
	 285.46 415.67 l
cp p3
np
  288.18 416.16 m
	 291.29 420.67 l
	 291.57 425.29 l
	 288.50 420.34 l
cp p3
np
  291.29 420.67 m
	 294.44 425.33 l
	 294.67 430.47 l
	 291.57 425.29 l
cp p3
np
  294.44 425.33 m
	 297.62 430.06 l
	 297.81 435.78 l
	 294.67 430.47 l
cp p3
np
  297.62 430.06 m
	 300.84 434.72 l
	 300.99 441.10 l
	 297.81 435.78 l
cp p3
np
  300.84 434.72 m
	 304.11 439.16 l
	 304.21 446.26 l
	 300.99 441.10 l
cp p3
np
  304.11 439.16 m
	 307.41 443.15 l
	 307.48 451.00 l
	 304.21 446.26 l
cp p3
np
  307.41 443.15 m
	 310.76 446.48 l
	 310.80 455.03 l
	 307.48 451.00 l
cp p3
np
  310.76 446.48 m
	 314.13 448.88 l
	 314.16 458.00 l
	 310.80 455.03 l
cp p3
np
  314.13 448.88 m
	 317.53 450.15 l
	 317.54 459.59 l
	 314.16 458.00 l
cp p3
np
  257.64 388.86 m
	 260.72 389.98 l
	 261.47 392.00 l
	 258.44 390.80 l
cp p3
np
  260.72 389.98 m
	 263.78 391.35 l
	 264.49 393.48 l
	 261.47 392.00 l
cp p3
np
  263.78 391.35 m
	 266.84 393.04 l
	 267.50 395.32 l
	 264.49 393.48 l
cp p3
np
  324.37 440.10 m
	 327.77 438.13 l
	 327.72 446.48 l
	 324.34 448.88 l
cp p3
np
  314.11 440.10 m
	 317.53 441.12 l
	 317.53 450.15 l
	 314.13 448.88 l
cp p3
np
  317.53 441.12 m
	 320.95 441.12 l
	 320.94 450.15 l
	 317.53 450.15 l
cp p3
np
  320.95 441.12 m
	 324.37 440.10 l
	 324.34 448.88 l
	 320.94 450.15 l
cp p3
np
  337.78 428.18 m
	 341.04 424.12 l
	 340.86 430.06 l
	 337.63 434.72 l
cp p3
np
  327.77 438.13 m
	 331.14 435.36 l
	 331.06 443.15 l
	 327.72 446.48 l
cp p3
np
  331.14 435.36 m
	 334.48 431.99 l
	 334.37 439.16 l
	 331.06 443.15 l
cp p3
np
  334.48 431.99 m
	 337.78 428.18 l
	 337.63 434.72 l
	 334.37 439.16 l
cp p3
np
  350.62 411.72 m
	 353.75 407.82 l
	 353.38 411.87 l
	 350.30 416.16 l
cp p3
np
  353.75 407.82 m
	 356.87 404.16 l
	 356.45 407.85 l
	 353.38 411.87 l
cp p3
np
  356.87 404.16 m
	 359.96 400.76 l
	 359.50 404.15 l
	 356.45 407.85 l
cp p3
np
  359.96 400.76 m
	 363.05 397.67 l
	 362.53 400.78 l
	 359.50 404.15 l
cp p3
np
  363.05 397.67 m
	 366.13 394.88 l
	 365.56 397.77 l
	 362.53 400.78 l
cp p3
np
  366.13 394.88 m
	 369.21 392.55 l
	 368.59 395.14 l
	 365.56 397.77 l
cp p3
np
  369.21 392.55 m
	 372.31 390.67 l
	 371.64 393.04 l
	 368.59 395.14 l
cp p3
np
  372.31 390.67 m
	 375.41 389.14 l
	 374.69 391.35 l
	 371.64 393.04 l
cp p3
np
  375.41 389.14 m
	 378.53 387.89 l
	 377.76 389.98 l
	 374.69 391.35 l
cp p3
np
  378.53 387.89 m
	 381.65 386.85 l
	 380.83 388.86 l
	 377.76 389.98 l
cp p3
np
  341.04 424.12 m
	 344.27 419.95 l
	 344.04 425.33 l
	 340.86 430.06 l
cp p3
np
  344.27 419.95 m
	 347.46 415.78 l
	 347.18 420.67 l
	 344.04 425.33 l
cp p3
np
  347.46 415.78 m
	 350.62 411.72 l
	 350.30 416.16 l
	 347.18 420.67 l
cp p3
np
  259.95 387.89 m
	 263.06 389.14 l
	 263.78 391.35 l
	 260.72 389.98 l
cp p3
np
  263.06 389.14 m
	 266.17 390.67 l
	 266.84 393.04 l
	 263.78 391.35 l
cp p3
np
  266.17 390.67 m
	 269.26 392.55 l
	 269.88 395.14 l
	 266.84 393.04 l
cp p3
np
  269.26 392.55 m
	 272.35 394.88 l
	 272.91 397.77 l
	 269.88 395.14 l
cp p3
np
  272.35 394.88 m
	 275.43 397.67 l
	 275.94 400.78 l
	 272.91 397.77 l
cp p3
np
  275.43 397.67 m
	 278.51 400.76 l
	 278.98 404.15 l
	 275.94 400.78 l
cp p3
np
  278.51 400.76 m
	 281.61 404.16 l
	 282.03 407.85 l
	 278.98 404.15 l
cp p3
np
  281.61 404.16 m
	 284.72 407.82 l
	 285.09 411.87 l
	 282.03 407.85 l
cp p3
np
  284.72 407.82 m
	 287.86 411.72 l
	 288.18 416.16 l
	 285.09 411.87 l
cp p3
np
  287.86 411.72 m
	 291.02 415.78 l
	 291.29 420.67 l
	 288.18 416.16 l
cp p3
np
  291.02 415.78 m
	 294.21 419.95 l
	 294.44 425.33 l
	 291.29 420.67 l
cp p3
np
  294.21 419.95 m
	 297.44 424.12 l
	 297.62 430.06 l
	 294.44 425.33 l
cp p3
np
  297.44 424.12 m
	 300.70 428.18 l
	 300.84 434.72 l
	 297.62 430.06 l
cp p3
np
  300.70 428.18 m
	 304.00 431.99 l
	 304.11 439.16 l
	 300.84 434.72 l
cp p3
np
  304.00 431.99 m
	 307.34 435.36 l
	 307.41 443.15 l
	 304.11 439.16 l
cp p3
np
  307.34 435.36 m
	 310.71 438.13 l
	 310.76 446.48 l
	 307.41 443.15 l
cp p3
np
  310.71 438.13 m
	 314.11 440.10 l
	 314.13 448.88 l
	 310.76 446.48 l
cp p3
np
  256.83 386.85 m
	 259.95 387.89 l
	 260.72 389.98 l
	 257.64 388.86 l
cp p3
np
  310.65 430.04 m
	 314.08 431.67 l
	 314.11 440.10 l
	 310.71 438.13 l
cp p3
np
  317.52 432.51 m
	 320.96 432.51 l
	 320.95 441.12 l
	 317.53 441.12 l
cp p3
np
  320.96 432.51 m
	 324.40 431.67 l
	 324.37 440.10 l
	 320.95 441.12 l
cp p3
np
  324.40 431.67 m
	 327.82 430.04 l
	 327.77 438.13 l
	 324.37 440.10 l
cp p3
np
  314.08 431.67 m
	 317.52 432.51 l
	 317.53 441.12 l
	 314.11 440.10 l
cp p3
np
  331.22 427.73 m
	 334.59 424.87 l
	 334.48 431.99 l
	 331.14 435.36 l
cp p3
np
  334.59 424.87 m
	 337.93 421.61 l
	 337.78 428.18 l
	 334.48 431.99 l
cp p3
np
  337.93 421.61 m
	 341.23 418.09 l
	 341.04 424.12 l
	 337.78 428.18 l
cp p3
np
  327.82 430.04 m
	 331.22 427.73 l
	 331.14 435.36 l
	 327.77 438.13 l
cp p3
np
  344.50 414.43 m
	 347.73 410.74 l
	 347.46 415.78 l
	 344.27 419.95 l
cp p3
np
  347.73 410.74 m
	 350.94 407.11 l
	 350.62 411.72 l
	 347.46 415.78 l
cp p3
np
  350.94 407.11 m
	 354.13 403.61 l
	 353.75 407.82 l
	 350.62 411.72 l
cp p3
np
  354.13 403.61 m
	 357.29 400.30 l
	 356.87 404.16 l
	 353.75 407.82 l
cp p3
np
  357.29 400.30 m
	 360.44 397.23 l
	 359.96 400.76 l
	 356.87 404.16 l
cp p3
np
  360.44 397.23 m
	 363.57 394.42 l
	 363.05 397.67 l
	 359.96 400.76 l
cp p3
np
  363.57 394.42 m
	 366.71 391.93 l
	 366.13 394.88 l
	 363.05 397.67 l
cp p3
np
  366.71 391.93 m
	 369.85 389.90 l
	 369.21 392.55 l
	 366.13 394.88 l
cp p3
np
  369.85 389.90 m
	 373.00 388.23 l
	 372.31 390.67 l
	 369.21 392.55 l
cp p3
np
  373.00 388.23 m
	 376.16 386.86 l
	 375.41 389.14 l
	 372.31 390.67 l
cp p3
np
  376.16 386.86 m
	 379.32 385.72 l
	 378.53 387.89 l
	 375.41 389.14 l
cp p3
np
  379.32 385.72 m
	 382.49 384.76 l
	 381.65 386.85 l
	 378.53 387.89 l
cp p3
np
  341.23 418.09 m
	 344.50 414.43 l
	 344.27 419.95 l
	 341.04 424.12 l
cp p3
np
  255.99 384.76 m
	 259.16 385.72 l
	 259.95 387.89 l
	 256.83 386.85 l
cp p3
np
  259.16 385.72 m
	 262.32 386.86 l
	 263.06 389.14 l
	 259.95 387.89 l
cp p3
np
  262.32 386.86 m
	 265.48 388.23 l
	 266.17 390.67 l
	 263.06 389.14 l
cp p3
np
  265.48 388.23 m
	 268.63 389.90 l
	 269.26 392.55 l
	 266.17 390.67 l
cp p3
np
  268.63 389.90 m
	 271.77 391.93 l
	 272.35 394.88 l
	 269.26 392.55 l
cp p3
np
  271.77 391.93 m
	 274.90 394.42 l
	 275.43 397.67 l
	 272.35 394.88 l
cp p3
np
  274.90 394.42 m
	 278.04 397.23 l
	 278.51 400.76 l
	 275.43 397.67 l
cp p3
np
  278.04 397.23 m
	 281.19 400.30 l
	 281.61 404.16 l
	 278.51 400.76 l
cp p3
np
  281.19 400.30 m
	 284.35 403.61 l
	 284.72 407.82 l
	 281.61 404.16 l
cp p3
np
  284.35 403.61 m
	 287.53 407.11 l
	 287.86 411.72 l
	 284.72 407.82 l
cp p3
np
  287.53 407.11 m
	 290.74 410.74 l
	 291.02 415.78 l
	 287.86 411.72 l
cp p3
np
  290.74 410.74 m
	 293.98 414.43 l
	 294.21 419.95 l
	 291.02 415.78 l
cp p3
np
  293.98 414.43 m
	 297.25 418.09 l
	 297.44 424.12 l
	 294.21 419.95 l
cp p3
np
  297.25 418.09 m
	 300.55 421.61 l
	 300.70 428.18 l
	 297.44 424.12 l
cp p3
np
  300.55 421.61 m
	 303.89 424.87 l
	 304.00 431.99 l
	 300.70 428.18 l
cp p3
np
  303.89 424.87 m
	 307.26 427.73 l
	 307.34 435.36 l
	 304.00 431.99 l
cp p3
np
  307.26 427.73 m
	 310.65 430.04 l
	 310.71 438.13 l
	 307.34 435.36 l
cp p3
np
  300.39 415.10 m
	 303.77 417.89 l
	 303.89 424.87 l
	 300.55 421.61 l
cp p3
np
  303.77 417.89 m
	 307.17 420.31 l
	 307.26 427.73 l
	 303.89 424.87 l
cp p3
np
  307.17 420.31 m
	 310.60 422.25 l
	 310.65 430.04 l
	 307.26 427.73 l
cp p3
np
  310.60 422.25 m
	 314.04 423.61 l
	 314.08 431.67 l
	 310.65 430.04 l
cp p3
np
  314.04 423.61 m
	 317.51 424.31 l
	 317.52 432.51 l
	 314.08 431.67 l
cp p3
np
  317.51 424.31 m
	 320.97 424.31 l
	 320.96 432.51 l
	 317.52 432.51 l
cp p3
np
  320.97 424.31 m
	 324.43 423.61 l
	 324.40 431.67 l
	 320.96 432.51 l
cp p3
np
  324.43 423.61 m
	 327.88 422.25 l
	 327.82 430.04 l
	 324.40 431.67 l
cp p3
np
  327.88 422.25 m
	 331.31 420.31 l
	 331.22 427.73 l
	 327.82 430.04 l
cp p3
np
  331.31 420.31 m
	 334.71 417.89 l
	 334.59 424.87 l
	 331.22 427.73 l
cp p3
np
  334.71 417.89 m
	 338.08 415.10 l
	 337.93 421.61 l
	 334.59 424.87 l
cp p3
np
  338.08 415.10 m
	 341.42 412.05 l
	 341.23 418.09 l
	 337.93 421.61 l
cp p3
np
  341.42 412.05 m
	 344.74 408.86 l
	 344.50 414.43 l
	 341.23 418.09 l
cp p3
np
  344.74 408.86 m
	 348.02 405.62 l
	 347.73 410.74 l
	 344.50 414.43 l
cp p3
np
  348.02 405.62 m
	 351.27 402.41 l
	 350.94 407.11 l
	 347.73 410.74 l
cp p3
np
  351.27 402.41 m
	 354.51 399.30 l
	 354.13 403.61 l
	 350.94 407.11 l
cp p3
np
  354.51 399.30 m
	 357.72 396.35 l
	 357.29 400.30 l
	 354.13 403.61 l
cp p3
np
  357.72 396.35 m
	 360.92 393.59 l
	 360.44 397.23 l
	 357.29 400.30 l
cp p3
np
  360.92 393.59 m
	 364.11 391.08 l
	 363.57 394.42 l
	 360.44 397.23 l
cp p3
np
  364.11 391.08 m
	 367.30 388.95 l
	 366.71 391.93 l
	 363.57 394.42 l
cp p3
np
  367.30 388.95 m
	 370.50 387.19 l
	 369.85 389.90 l
	 366.71 391.93 l
cp p3
np
  370.50 387.19 m
	 373.71 385.73 l
	 373.00 388.23 l
	 369.85 389.90 l
cp p3
np
  373.71 385.73 m
	 376.92 384.51 l
	 376.16 386.86 l
	 373.00 388.23 l
cp p3
np
  376.92 384.51 m
	 380.13 383.48 l
	 379.32 385.72 l
	 376.16 386.86 l
cp p3
np
  380.13 383.48 m
	 383.35 382.62 l
	 382.49 384.76 l
	 379.32 385.72 l
cp p3
np
  293.74 408.86 m
	 297.05 412.05 l
	 297.25 418.09 l
	 293.98 414.43 l
cp p3
np
  255.12 382.62 m
	 258.34 383.48 l
	 259.16 385.72 l
	 255.99 384.76 l
cp p3
np
  258.34 383.48 m
	 261.56 384.51 l
	 262.32 386.86 l
	 259.16 385.72 l
cp p3
np
  261.56 384.51 m
	 264.77 385.73 l
	 265.48 388.23 l
	 262.32 386.86 l
cp p3
np
  264.77 385.73 m
	 267.97 387.19 l
	 268.63 389.90 l
	 265.48 388.23 l
cp p3
np
  267.97 387.19 m
	 271.17 388.95 l
	 271.77 391.93 l
	 268.63 389.90 l
cp p3
np
  271.17 388.95 m
	 274.36 391.08 l
	 274.90 394.42 l
	 271.77 391.93 l
cp p3
np
  274.36 391.08 m
	 277.55 393.59 l
	 278.04 397.23 l
	 274.90 394.42 l
cp p3
np
  277.55 393.59 m
	 280.75 396.35 l
	 281.19 400.30 l
	 278.04 397.23 l
cp p3
np
  280.75 396.35 m
	 283.97 399.30 l
	 284.35 403.61 l
	 281.19 400.30 l
cp p3
np
  283.97 399.30 m
	 287.20 402.41 l
	 287.53 407.11 l
	 284.35 403.61 l
cp p3
np
  287.20 402.41 m
	 290.46 405.62 l
	 290.74 410.74 l
	 287.53 407.11 l
cp p3
np
  290.46 405.62 m
	 293.74 408.86 l
	 293.98 414.43 l
	 290.74 410.74 l
cp p3
np
  297.05 412.05 m
	 300.39 415.10 l
	 300.55 421.61 l
	 297.25 418.09 l
cp p3
np
  380.97 381.19 m
	 384.24 380.41 l
	 383.35 382.62 l
	 380.13 383.48 l
cp p3
np
  296.85 406.10 m
	 300.23 408.71 l
	 300.39 415.10 l
	 297.05 412.05 l
cp p3
np
  300.23 408.71 m
	 303.64 411.10 l
	 303.77 417.89 l
	 300.39 415.10 l
cp p3
np
  303.64 411.10 m
	 307.08 413.15 l
	 307.17 420.31 l
	 303.77 417.89 l
cp p3
np
  307.08 413.15 m
	 310.53 414.79 l
	 310.60 422.25 l
	 307.17 420.31 l
cp p3
np
  310.53 414.79 m
	 314.01 415.93 l
	 314.04 423.61 l
	 310.60 422.25 l
cp p3
np
  314.01 415.93 m
	 317.49 416.51 l
	 317.51 424.31 l
	 314.04 423.61 l
cp p3
np
  317.49 416.51 m
	 320.98 416.51 l
	 320.97 424.31 l
	 317.51 424.31 l
cp p3
np
  320.98 416.51 m
	 324.47 415.93 l
	 324.43 423.61 l
	 320.97 424.31 l
cp p3
np
  324.47 415.93 m
	 327.94 414.79 l
	 327.88 422.25 l
	 324.43 423.61 l
cp p3
np
  327.94 414.79 m
	 331.40 413.15 l
	 331.31 420.31 l
	 327.88 422.25 l
cp p3
np
  331.40 413.15 m
	 334.84 411.10 l
	 334.71 417.89 l
	 331.31 420.31 l
cp p3
np
  334.84 411.10 m
	 338.24 408.71 l
	 338.08 415.10 l
	 334.71 417.89 l
cp p3
np
  338.24 408.71 m
	 341.63 406.10 l
	 341.42 412.05 l
	 338.08 415.10 l
cp p3
np
  341.63 406.10 m
	 344.98 403.33 l
	 344.74 408.86 l
	 341.42 412.05 l
cp p3
np
  344.98 403.33 m
	 348.31 400.50 l
	 348.02 405.62 l
	 344.74 408.86 l
cp p3
np
  348.31 400.50 m
	 351.62 397.69 l
	 351.27 402.41 l
	 348.02 405.62 l
cp p3
np
  351.62 397.69 m
	 354.90 394.95 l
	 354.51 399.30 l
	 351.27 402.41 l
cp p3
np
  354.90 394.95 m
	 358.17 392.34 l
	 357.72 396.35 l
	 354.51 399.30 l
cp p3
np
  358.17 392.34 m
	 361.42 389.90 l
	 360.92 393.59 l
	 357.72 396.35 l
cp p3
np
  361.42 389.90 m
	 364.67 387.77 l
	 364.11 391.08 l
	 360.92 393.59 l
cp p3
np
  364.67 387.77 m
	 367.92 385.98 l
	 367.30 388.95 l
	 364.11 391.08 l
cp p3
np
  367.92 385.98 m
	 371.18 384.46 l
	 370.50 387.19 l
	 367.30 388.95 l
cp p3
np
  371.18 384.46 m
	 374.44 383.19 l
	 373.71 385.73 l
	 370.50 387.19 l
cp p3
np
  374.44 383.19 m
	 377.70 382.11 l
	 376.92 384.51 l
	 373.71 385.73 l
cp p3
np
  377.70 382.11 m
	 380.97 381.19 l
	 380.13 383.48 l
	 376.92 384.51 l
cp p3
np
  283.58 394.95 m
	 286.86 397.69 l
	 287.20 402.41 l
	 283.97 399.30 l
cp p3
np
  286.86 397.69 m
	 290.17 400.50 l
	 290.46 405.62 l
	 287.20 402.41 l
cp p3
np
  290.17 400.50 m
	 293.49 403.33 l
	 293.74 408.86 l
	 290.46 405.62 l
cp p3
np
  293.49 403.33 m
	 296.85 406.10 l
	 297.05 412.05 l
	 293.74 408.86 l
cp p3
np
  254.24 380.41 m
	 257.51 381.19 l
	 258.34 383.48 l
	 255.12 382.62 l
cp p3
np
  257.51 381.19 m
	 260.78 382.11 l
	 261.56 384.51 l
	 258.34 383.48 l
cp p3
np
  260.78 382.11 m
	 264.04 383.19 l
	 264.77 385.73 l
	 261.56 384.51 l
cp p3
np
  264.04 383.19 m
	 267.30 384.46 l
	 267.97 387.19 l
	 264.77 385.73 l
cp p3
np
  267.30 384.46 m
	 270.55 385.98 l
	 271.17 388.95 l
	 267.97 387.19 l
cp p3
np
  270.55 385.98 m
	 273.81 387.77 l
	 274.36 391.08 l
	 271.17 388.95 l
cp p3
np
  273.81 387.77 m
	 277.06 389.90 l
	 277.55 393.59 l
	 274.36 391.08 l
cp p3
np
  277.06 389.90 m
	 280.31 392.34 l
	 280.75 396.35 l
	 277.55 393.59 l
cp p3
np
  280.31 392.34 m
	 283.58 394.95 l
	 283.97 399.30 l
	 280.75 396.35 l
cp p3
np
  371.87 381.72 m
	 375.19 380.61 l
	 374.44 383.19 l
	 371.18 384.46 l
cp p3
np
  375.19 380.61 m
	 378.51 379.66 l
	 377.70 382.11 l
	 374.44 383.19 l
cp p3
np
  378.51 379.66 m
	 381.83 378.85 l
	 380.97 381.19 l
	 377.70 382.11 l
cp p3
np
  381.83 378.85 m
	 385.15 378.15 l
	 384.24 380.41 l
	 380.97 381.19 l
cp p3
np
  293.24 397.89 m
	 296.63 400.27 l
	 296.85 406.10 l
	 293.49 403.33 l
cp p3
np
  296.63 400.27 m
	 300.06 402.51 l
	 300.23 408.71 l
	 296.85 406.10 l
cp p3
np
  300.06 402.51 m
	 303.50 404.54 l
	 303.64 411.10 l
	 300.23 408.71 l
cp p3
np
  303.50 404.54 m
	 306.97 406.28 l
	 307.08 413.15 l
	 303.64 411.10 l
cp p3
np
  306.97 406.28 m
	 310.46 407.66 l
	 310.53 414.79 l
	 307.08 413.15 l
cp p3
np
  310.46 407.66 m
	 313.97 408.62 l
	 314.01 415.93 l
	 310.53 414.79 l
cp p3
np
  313.97 408.62 m
	 317.48 409.11 l
	 317.49 416.51 l
	 314.01 415.93 l
cp p3
np
  317.48 409.11 m
	 321.00 409.11 l
	 320.98 416.51 l
	 317.49 416.51 l
cp p3
np
  321.00 409.11 m
	 324.51 408.62 l
	 324.47 415.93 l
	 320.98 416.51 l
cp p3
np
  324.51 408.62 m
	 328.01 407.66 l
	 327.94 414.79 l
	 324.47 415.93 l
cp p3
np
  328.01 407.66 m
	 331.50 406.28 l
	 331.40 413.15 l
	 327.94 414.79 l
cp p3
np
  331.50 406.28 m
	 334.97 404.54 l
	 334.84 411.10 l
	 331.40 413.15 l
cp p3
np
  334.97 404.54 m
	 338.42 402.51 l
	 338.24 408.71 l
	 334.84 411.10 l
cp p3
np
  338.42 402.51 m
	 341.84 400.27 l
	 341.63 406.10 l
	 338.24 408.71 l
cp p3
np
  341.84 400.27 m
	 345.24 397.89 l
	 344.98 403.33 l
	 341.63 406.10 l
cp p3
np
  345.24 397.89 m
	 348.62 395.44 l
	 348.31 400.50 l
	 344.98 403.33 l
cp p3
np
  348.62 395.44 m
	 351.97 393.00 l
	 351.62 397.69 l
	 348.31 400.50 l
cp p3
np
  351.97 393.00 m
	 355.30 390.61 l
	 354.90 394.95 l
	 351.62 397.69 l
cp p3
np
  355.30 390.61 m
	 358.62 388.33 l
	 358.17 392.34 l
	 354.90 394.95 l
cp p3
np
  358.62 388.33 m
	 361.94 386.29 l
	 361.42 389.90 l
	 358.17 392.34 l
cp p3
np
  361.94 386.29 m
	 365.25 384.52 l
	 364.67 387.77 l
	 361.42 389.90 l
cp p3
np
  365.25 384.52 m
	 368.56 383.01 l
	 367.92 385.98 l
	 364.67 387.77 l
cp p3
np
  368.56 383.01 m
	 371.87 381.72 l
	 371.18 384.46 l
	 367.92 385.98 l
cp p3
np
  279.85 388.33 m
	 283.17 390.61 l
	 283.58 394.95 l
	 280.31 392.34 l
cp p3
np
  283.17 390.61 m
	 286.51 393.00 l
	 286.86 397.69 l
	 283.58 394.95 l
cp p3
np
  286.51 393.00 m
	 289.86 395.44 l
	 290.17 400.50 l
	 286.86 397.69 l
cp p3
np
  289.86 395.44 m
	 293.24 397.89 l
	 293.49 403.33 l
	 290.17 400.50 l
cp p3
np
  263.29 380.61 m
	 266.60 381.72 l
	 267.30 384.46 l
	 264.04 383.19 l
cp p3
np
  253.33 378.15 m
	 256.65 378.85 l
	 257.51 381.19 l
	 254.24 380.41 l
cp p3
np
  256.65 378.85 m
	 259.97 379.66 l
	 260.78 382.11 l
	 257.51 381.19 l
cp p3
np
  259.97 379.66 m
	 263.29 380.61 l
	 264.04 383.19 l
	 260.78 382.11 l
cp p3
np
  276.54 386.29 m
	 279.85 388.33 l
	 280.31 392.34 l
	 277.06 389.90 l
cp p3
np
  266.60 381.72 m
	 269.92 383.01 l
	 270.55 385.98 l
	 267.30 384.46 l
cp p3
np
  269.92 383.01 m
	 273.23 384.52 l
	 273.81 387.77 l
	 270.55 385.98 l
cp p3
np
  273.23 384.52 m
	 276.54 386.29 l
	 277.06 389.90 l
	 273.81 387.77 l
cp p3
np
  382.71 376.46 m
	 386.09 375.83 l
	 385.15 378.15 l
	 381.83 378.85 l
cp p3
np
  369.22 380.07 m
	 372.59 378.97 l
	 371.87 381.72 l
	 368.56 383.01 l
cp p3
np
  372.59 378.97 m
	 375.96 378.01 l
	 375.19 380.61 l
	 371.87 381.72 l
cp p3
np
  375.96 378.01 m
	 379.34 377.18 l
	 378.51 379.66 l
	 375.19 380.61 l
cp p3
np
  379.34 377.18 m
	 382.71 376.46 l
	 381.83 378.85 l
	 378.51 379.66 l
cp p3
np
  286.14 388.39 m
	 289.54 390.49 l
	 289.86 395.44 l
	 286.51 393.00 l
cp p3
np
  289.54 390.49 m
	 292.96 392.59 l
	 293.24 397.89 l
	 289.86 395.44 l
cp p3
np
  292.96 392.59 m
	 296.41 394.62 l
	 296.63 400.27 l
	 293.24 397.89 l
cp p3
np
  296.41 394.62 m
	 299.87 396.53 l
	 300.06 402.51 l
	 296.63 400.27 l
cp p3
np
  299.87 396.53 m
	 303.36 398.25 l
	 303.50 404.54 l
	 300.06 402.51 l
cp p3
np
  303.36 398.25 m
	 306.86 399.73 l
	 306.97 406.28 l
	 303.50 404.54 l
cp p3
np
  306.86 399.73 m
	 310.39 400.89 l
	 310.46 407.66 l
	 306.97 406.28 l
cp p3
np
  310.39 400.89 m
	 313.92 401.69 l
	 313.97 408.62 l
	 310.46 407.66 l
cp p3
np
  313.92 401.69 m
	 317.46 402.10 l
	 317.48 409.11 l
	 313.97 408.62 l
cp p3
np
  317.46 402.10 m
	 321.01 402.10 l
	 321.00 409.11 l
	 317.48 409.11 l
cp p3
np
  321.01 402.10 m
	 324.55 401.69 l
	 324.51 408.62 l
	 321.00 409.11 l
cp p3
np
  324.55 401.69 m
	 328.09 400.89 l
	 328.01 407.66 l
	 324.51 408.62 l
cp p3
np
  328.09 400.89 m
	 331.61 399.73 l
	 331.50 406.28 l
	 328.01 407.66 l
cp p3
np
  331.61 399.73 m
	 335.12 398.25 l
	 334.97 404.54 l
	 331.50 406.28 l
cp p3
np
  335.12 398.25 m
	 338.60 396.53 l
	 338.42 402.51 l
	 334.97 404.54 l
cp p3
np
  338.60 396.53 m
	 342.07 394.62 l
	 341.84 400.27 l
	 338.42 402.51 l
cp p3
np
  342.07 394.62 m
	 345.51 392.59 l
	 345.24 397.89 l
	 341.84 400.27 l
cp p3
np
  345.51 392.59 m
	 348.94 390.49 l
	 348.62 395.44 l
	 345.24 397.89 l
cp p3
np
  348.94 390.49 m
	 352.34 388.39 l
	 351.97 393.00 l
	 348.62 395.44 l
cp p3
np
  352.34 388.39 m
	 355.73 386.33 l
	 355.30 390.61 l
	 351.97 393.00 l
cp p3
np
  355.73 386.33 m
	 359.11 384.45 l
	 358.62 388.33 l
	 355.30 390.61 l
cp p3
np
  359.11 384.45 m
	 362.48 382.79 l
	 361.94 386.29 l
	 358.62 388.33 l
cp p3
np
  362.48 382.79 m
	 365.85 381.34 l
	 365.25 384.52 l
	 361.94 386.29 l
cp p3
np
  365.85 381.34 m
	 369.22 380.07 l
	 368.56 383.01 l
	 365.25 384.52 l
cp p3
np
  276.00 382.79 m
	 279.37 384.45 l
	 279.85 388.33 l
	 276.54 386.29 l
cp p3
np
  279.37 384.45 m
	 282.75 386.33 l
	 283.17 390.61 l
	 279.85 388.33 l
cp p3
np
  282.75 386.33 m
	 286.14 388.39 l
	 286.51 393.00 l
	 283.17 390.61 l
cp p3
np
  255.76 376.46 m
	 259.14 377.18 l
	 259.97 379.66 l
	 256.65 378.85 l
cp p3
np
  259.14 377.18 m
	 262.51 378.01 l
	 263.29 380.61 l
	 259.97 379.66 l
cp p3
np
  262.51 378.01 m
	 265.88 378.97 l
	 266.60 381.72 l
	 263.29 380.61 l
cp p3
np
  252.39 375.83 m
	 255.76 376.46 l
	 256.65 378.85 l
	 253.33 378.15 l
cp p3
np
  269.25 380.07 m
	 272.62 381.34 l
	 273.23 384.52 l
	 269.92 383.01 l
cp p3
np
  272.62 381.34 m
	 276.00 382.79 l
	 276.54 386.29 l
	 273.23 384.52 l
cp p3
np
  265.88 378.97 m
	 269.25 380.07 l
	 269.92 383.01 l
	 266.60 381.72 l
cp p3
np
  383.62 374.02 m
	 387.05 373.47 l
	 386.09 375.83 l
	 382.71 376.46 l
cp p3
np
  376.77 375.38 m
	 380.19 374.66 l
	 379.34 377.18 l
	 375.96 378.01 l
cp p3
np
  380.19 374.66 m
	 383.62 374.02 l
	 382.71 376.46 l
	 379.34 377.18 l
cp p3
np
  366.48 378.21 m
	 369.91 377.14 l
	 369.22 380.07 l
	 365.85 381.34 l
cp p3
np
  369.91 377.14 m
	 373.34 376.21 l
	 372.59 378.97 l
	 369.22 380.07 l
cp p3
np
  373.34 376.21 m
	 376.77 375.38 l
	 375.96 378.01 l
	 372.59 378.97 l
cp p3
np
  282.30 382.26 m
	 285.75 383.91 l
	 286.14 388.39 l
	 282.75 386.33 l
cp p3
np
  285.75 383.91 m
	 289.20 385.69 l
	 289.54 390.49 l
	 286.14 388.39 l
cp p3
np
  289.20 385.69 m
	 292.68 387.46 l
	 292.96 392.59 l
	 289.54 390.49 l
cp p3
np
  292.68 387.46 m
	 296.17 389.19 l
	 296.41 394.62 l
	 292.96 392.59 l
cp p3
np
  296.17 389.19 m
	 299.68 390.80 l
	 299.87 396.53 l
	 296.41 394.62 l
cp p3
np
  299.68 390.80 m
	 303.20 392.25 l
	 303.36 398.25 l
	 299.87 396.53 l
cp p3
np
  303.20 392.25 m
	 306.75 393.49 l
	 306.86 399.73 l
	 303.36 398.25 l
cp p3
np
  306.75 393.49 m
	 310.30 394.46 l
	 310.39 400.89 l
	 306.86 399.73 l
cp p3
np
  310.30 394.46 m
	 313.87 395.14 l
	 313.92 401.69 l
	 310.39 400.89 l
cp p3
np
  313.87 395.14 m
	 317.45 395.48 l
	 317.46 402.10 l
	 313.92 401.69 l
cp p3
np
  317.45 395.48 m
	 321.03 395.48 l
	 321.01 402.10 l
	 317.46 402.10 l
cp p3
np
  321.03 395.48 m
	 324.60 395.14 l
	 324.55 401.69 l
	 321.01 402.10 l
cp p3
np
  324.60 395.14 m
	 328.17 394.46 l
	 328.09 400.89 l
	 324.55 401.69 l
cp p3
np
  328.17 394.46 m
	 331.73 393.49 l
	 331.61 399.73 l
	 328.09 400.89 l
cp p3
np
  331.73 393.49 m
	 335.27 392.25 l
	 335.12 398.25 l
	 331.61 399.73 l
cp p3
np
  335.27 392.25 m
	 338.80 390.80 l
	 338.60 396.53 l
	 335.12 398.25 l
cp p3
np
  338.80 390.80 m
	 342.31 389.19 l
	 342.07 394.62 l
	 338.60 396.53 l
cp p3
np
  342.31 389.19 m
	 345.80 387.46 l
	 345.51 392.59 l
	 342.07 394.62 l
cp p3
np
  345.80 387.46 m
	 349.27 385.69 l
	 348.94 390.49 l
	 345.51 392.59 l
cp p3
np
  349.27 385.69 m
	 352.73 383.91 l
	 352.34 388.39 l
	 348.94 390.49 l
cp p3
np
  352.73 383.91 m
	 356.18 382.26 l
	 355.73 386.33 l
	 352.34 388.39 l
cp p3
np
  356.18 382.26 m
	 359.61 380.76 l
	 359.11 384.45 l
	 355.73 386.33 l
cp p3
np
  359.61 380.76 m
	 363.05 379.41 l
	 362.48 382.79 l
	 359.11 384.45 l
cp p3
np
  363.05 379.41 m
	 366.48 378.21 l
	 365.85 381.34 l
	 362.48 382.79 l
cp p3
np
  268.57 377.14 m
	 272.00 378.21 l
	 272.62 381.34 l
	 269.25 380.07 l
cp p3
np
  272.00 378.21 m
	 275.43 379.41 l
	 276.00 382.79 l
	 272.62 381.34 l
cp p3
np
  275.43 379.41 m
	 278.86 380.76 l
	 279.37 384.45 l
	 276.00 382.79 l
cp p3
np
  278.86 380.76 m
	 282.30 382.26 l
	 282.75 386.33 l
	 279.37 384.45 l
cp p3
np
  251.42 373.47 m
	 254.85 374.02 l
	 255.76 376.46 l
	 252.39 375.83 l
cp p3
np
  254.85 374.02 m
	 258.28 374.66 l
	 259.14 377.18 l
	 255.76 376.46 l
cp p3
np
  258.28 374.66 m
	 261.71 375.38 l
	 262.51 378.01 l
	 259.14 377.18 l
cp p3
np
  261.71 375.38 m
	 265.14 376.21 l
	 265.88 378.97 l
	 262.51 378.01 l
cp p3
np
  265.14 376.21 m
	 268.57 377.14 l
	 269.25 380.07 l
	 265.88 378.97 l
cp p3
np
  377.59 372.73 m
	 381.08 372.10 l
	 380.19 374.66 l
	 376.77 375.38 l
cp p3
np
  381.08 372.10 m
	 384.56 371.54 l
	 383.62 374.02 l
	 380.19 374.66 l
cp p3
np
  384.56 371.54 m
	 388.05 371.05 l
	 387.05 373.47 l
	 383.62 374.02 l
cp p3
np
  374.11 373.44 m
	 377.59 372.73 l
	 376.77 375.38 l
	 373.34 376.21 l
cp p3
np
  360.15 377.22 m
	 363.64 376.12 l
	 363.05 379.41 l
	 359.61 380.76 l
cp p3
np
  363.64 376.12 m
	 367.13 375.13 l
	 366.48 378.21 l
	 363.05 379.41 l
cp p3
np
  367.13 375.13 m
	 370.62 374.24 l
	 369.91 377.14 l
	 366.48 378.21 l
cp p3
np
  370.62 374.24 m
	 374.11 373.44 l
	 373.34 376.21 l
	 369.91 377.14 l
cp p3
np
  278.33 377.22 m
	 281.83 378.42 l
	 282.30 382.26 l
	 278.86 380.76 l
cp p3
np
  281.83 378.42 m
	 285.33 379.72 l
	 285.75 383.91 l
	 282.30 382.26 l
cp p3
np
  285.33 379.72 m
	 288.85 381.10 l
	 289.20 385.69 l
	 285.75 383.91 l
cp p3
np
  288.85 381.10 m
	 292.37 382.55 l
	 292.68 387.46 l
	 289.20 385.69 l
cp p3
np
  292.37 382.55 m
	 295.91 384.00 l
	 296.17 389.19 l
	 292.68 387.46 l
cp p3
np
  295.91 384.00 m
	 299.46 385.34 l
	 299.68 390.80 l
	 296.17 389.19 l
cp p3
np
  299.46 385.34 m
	 303.03 386.56 l
	 303.20 392.25 l
	 299.68 390.80 l
cp p3
np
  303.03 386.56 m
	 306.62 387.59 l
	 306.75 393.49 l
	 303.20 392.25 l
cp p3
np
  306.62 387.59 m
	 310.21 388.40 l
	 310.30 394.46 l
	 306.75 393.49 l
cp p3
np
  310.21 388.40 m
	 313.82 388.96 l
	 313.87 395.14 l
	 310.30 394.46 l
cp p3
np
  313.82 388.96 m
	 317.43 389.25 l
	 317.45 395.48 l
	 313.87 395.14 l
cp p3
np
  317.43 389.25 m
	 321.04 389.25 l
	 321.03 395.48 l
	 317.45 395.48 l
cp p3
np
  321.04 389.25 m
	 324.66 388.96 l
	 324.60 395.14 l
	 321.03 395.48 l
cp p3
np
  324.66 388.96 m
	 328.26 388.40 l
	 328.17 394.46 l
	 324.60 395.14 l
cp p3
np
  328.26 388.40 m
	 331.86 387.59 l
	 331.73 393.49 l
	 328.17 394.46 l
cp p3
np
  331.86 387.59 m
	 335.44 386.56 l
	 335.27 392.25 l
	 331.73 393.49 l
cp p3
np
  335.44 386.56 m
	 339.01 385.34 l
	 338.80 390.80 l
	 335.27 392.25 l
cp p3
np
  339.01 385.34 m
	 342.57 384.00 l
	 342.31 389.19 l
	 338.80 390.80 l
cp p3
np
  342.57 384.00 m
	 346.10 382.55 l
	 345.80 387.46 l
	 342.31 389.19 l
cp p3
np
  346.10 382.55 m
	 349.63 381.10 l
	 349.27 385.69 l
	 345.80 387.46 l
cp p3
np
  349.63 381.10 m
	 353.14 379.72 l
	 352.73 383.91 l
	 349.27 385.69 l
cp p3
np
  353.14 379.72 m
	 356.65 378.42 l
	 356.18 382.26 l
	 352.73 383.91 l
cp p3
np
  356.65 378.42 m
	 360.15 377.22 l
	 359.61 380.76 l
	 356.18 382.26 l
cp p3
np
  264.37 373.44 m
	 267.85 374.24 l
	 268.57 377.14 l
	 265.14 376.21 l
cp p3
np
  267.85 374.24 m
	 271.34 375.13 l
	 272.00 378.21 l
	 268.57 377.14 l
cp p3
np
  271.34 375.13 m
	 274.83 376.12 l
	 275.43 379.41 l
	 272.00 378.21 l
cp p3
np
  274.83 376.12 m
	 278.33 377.22 l
	 278.86 380.76 l
	 275.43 379.41 l
cp p3
np
  260.88 372.73 m
	 264.37 373.44 l
	 265.14 376.21 l
	 261.71 375.38 l
cp p3
np
  250.42 371.05 m
	 253.91 371.54 l
	 254.85 374.02 l
	 251.42 373.47 l
cp p3
np
  253.91 371.54 m
	 257.40 372.10 l
	 258.28 374.66 l
	 254.85 374.02 l
cp p3
np
  257.40 372.10 m
	 260.88 372.73 l
	 261.71 375.38 l
	 258.28 374.66 l
cp p3
np
  371.36 371.34 m
	 374.91 370.66 l
	 374.11 373.44 l
	 370.62 374.24 l
cp p3
np
  374.91 370.66 m
	 378.45 370.05 l
	 377.59 372.73 l
	 374.11 373.44 l
cp p3
np
  378.45 370.05 m
	 381.99 369.51 l
	 381.08 372.10 l
	 377.59 372.73 l
cp p3
np
  381.99 369.51 m
	 385.54 369.02 l
	 384.56 371.54 l
	 381.08 372.10 l
cp p3
np
  385.54 369.02 m
	 389.08 368.58 l
	 388.05 371.05 l
	 384.56 371.54 l
cp p3
np
  357.15 374.77 m
	 360.71 373.81 l
	 360.15 377.22 l
	 356.65 378.42 l
cp p3
np
  360.71 373.81 m
	 364.26 372.91 l
	 363.64 376.12 l
	 360.15 377.22 l
cp p3
np
  364.26 372.91 m
	 367.81 372.09 l
	 367.13 375.13 l
	 363.64 376.12 l
cp p3
np
  367.81 372.09 m
	 371.36 371.34 l
	 370.62 374.24 l
	 367.13 375.13 l
cp p3
np
  270.66 372.09 m
	 274.21 372.91 l
	 274.83 376.12 l
	 271.34 375.13 l
cp p3
np
  274.21 372.91 m
	 277.77 373.81 l
	 278.33 377.22 l
	 274.83 376.12 l
cp p3
np
  277.77 373.81 m
	 281.32 374.77 l
	 281.83 378.42 l
	 278.33 377.22 l
cp p3
np
  281.32 374.77 m
	 284.89 375.80 l
	 285.33 379.72 l
	 281.83 378.42 l
cp p3
np
  284.89 375.80 m
	 288.46 376.88 l
	 288.85 381.10 l
	 285.33 379.72 l
cp p3
np
  288.46 376.88 m
	 292.04 377.99 l
	 292.37 382.55 l
	 288.85 381.10 l
cp p3
np
  292.04 377.99 m
	 295.63 379.10 l
	 295.91 384.00 l
	 292.37 382.55 l
cp p3
np
  295.63 379.10 m
	 299.24 380.18 l
	 299.46 385.34 l
	 295.91 384.00 l
cp p3
np
  299.24 380.18 m
	 302.85 381.18 l
	 303.03 386.56 l
	 299.46 385.34 l
cp p3
np
  302.85 381.18 m
	 306.48 382.03 l
	 306.62 387.59 l
	 303.03 386.56 l
cp p3
np
  306.48 382.03 m
	 310.12 382.70 l
	 310.21 388.40 l
	 306.62 387.59 l
cp p3
np
  310.12 382.70 m
	 313.76 383.16 l
	 313.82 388.96 l
	 310.21 388.40 l
cp p3
np
  313.76 383.16 m
	 317.41 383.40 l
	 317.43 389.25 l
	 313.82 388.96 l
cp p3
np
  317.41 383.40 m
	 321.06 383.40 l
	 321.04 389.25 l
	 317.43 389.25 l
cp p3
np
  321.06 383.40 m
	 324.71 383.16 l
	 324.66 388.96 l
	 321.04 389.25 l
cp p3
np
  324.71 383.16 m
	 328.36 382.70 l
	 328.26 388.40 l
	 324.66 388.96 l
cp p3
np
  328.36 382.70 m
	 332.00 382.03 l
	 331.86 387.59 l
	 328.26 388.40 l
cp p3
np
  332.00 382.03 m
	 335.62 381.18 l
	 335.44 386.56 l
	 331.86 387.59 l
cp p3
np
  335.62 381.18 m
	 339.24 380.18 l
	 339.01 385.34 l
	 335.44 386.56 l
cp p3
np
  339.24 380.18 m
	 342.84 379.10 l
	 342.57 384.00 l
	 339.01 385.34 l
cp p3
np
  342.84 379.10 m
	 346.43 377.99 l
	 346.10 382.55 l
	 342.57 384.00 l
cp p3
np
  346.43 377.99 m
	 350.01 376.88 l
	 349.63 381.10 l
	 346.10 382.55 l
cp p3
np
  350.01 376.88 m
	 353.59 375.80 l
	 353.14 379.72 l
	 349.63 381.10 l
cp p3
np
  353.59 375.80 m
	 357.15 374.77 l
	 356.65 378.42 l
	 353.14 379.72 l
cp p3
np
  260.03 370.05 m
	 263.57 370.66 l
	 264.37 373.44 l
	 260.88 372.73 l
cp p3
np
  263.57 370.66 m
	 267.12 371.34 l
	 267.85 374.24 l
	 264.37 373.44 l
cp p3
np
  267.12 371.34 m
	 270.66 372.09 l
	 271.34 375.13 l
	 267.85 374.24 l
cp p3
np
  252.94 369.02 m
	 256.48 369.51 l
	 257.40 372.10 l
	 253.91 371.54 l
cp p3
np
  256.48 369.51 m
	 260.03 370.05 l
	 260.88 372.73 l
	 257.40 372.10 l
cp p3
np
  249.40 368.58 m
	 252.94 369.02 l
	 253.91 371.54 l
	 250.42 371.05 l
cp p3
np
  372.13 368.45 m
	 375.73 367.87 l
	 374.91 370.66 l
	 371.36 371.34 l
cp p3
np
  364.91 369.76 m
	 368.52 369.08 l
	 367.81 372.09 l
	 364.26 372.91 l
cp p3
np
  368.52 369.08 m
	 372.13 368.45 l
	 371.36 371.34 l
	 367.81 372.09 l
cp p3
np
  386.54 366.45 m
	 390.14 366.06 l
	 389.08 368.58 l
	 385.54 369.02 l
cp p3
np
  375.73 367.87 m
	 379.34 367.35 l
	 378.45 370.05 l
	 374.91 370.66 l
cp p3
np
  379.34 367.35 m
	 382.94 366.87 l
	 381.99 369.51 l
	 378.45 370.05 l
cp p3
np
  382.94 366.87 m
	 386.54 366.45 l
	 385.54 369.02 l
	 381.99 369.51 l
cp p3
np
  354.06 372.10 m
	 357.68 371.27 l
	 357.15 374.77 l
	 353.59 375.80 l
cp p3
np
  357.68 371.27 m
	 361.30 370.49 l
	 360.71 373.81 l
	 357.15 374.77 l
cp p3
np
  361.30 370.49 m
	 364.91 369.76 l
	 364.26 372.91 l
	 360.71 373.81 l
cp p3
np
  266.35 368.45 m
	 269.95 369.08 l
	 270.66 372.09 l
	 267.12 371.34 l
cp p3
np
  269.95 369.08 m
	 273.56 369.76 l
	 274.21 372.91 l
	 270.66 372.09 l
cp p3
np
  273.56 369.76 m
	 277.18 370.49 l
	 277.77 373.81 l
	 274.21 372.91 l
cp p3
np
  277.18 370.49 m
	 280.80 371.27 l
	 281.32 374.77 l
	 277.77 373.81 l
cp p3
np
  280.80 371.27 m
	 284.42 372.10 l
	 284.89 375.80 l
	 281.32 374.77 l
cp p3
np
  284.42 372.10 m
	 288.05 372.95 l
	 288.46 376.88 l
	 284.89 375.80 l
cp p3
np
  288.05 372.95 m
	 291.69 373.81 l
	 292.04 377.99 l
	 288.46 376.88 l
cp p3
np
  291.69 373.81 m
	 295.33 374.66 l
	 295.63 379.10 l
	 292.04 377.99 l
cp p3
np
  295.33 374.66 m
	 298.99 375.47 l
	 299.24 380.18 l
	 295.63 379.10 l
cp p3
np
  298.99 375.47 m
	 302.66 376.22 l
	 302.85 381.18 l
	 299.24 380.18 l
cp p3
np
  302.66 376.22 m
	 306.33 376.87 l
	 306.48 382.03 l
	 302.85 381.18 l
cp p3
np
  306.33 376.87 m
	 310.01 377.38 l
	 310.12 382.70 l
	 306.48 382.03 l
cp p3
np
  310.01 377.38 m
	 313.70 377.75 l
	 313.76 383.16 l
	 310.12 382.70 l
cp p3
np
  313.70 377.75 m
	 317.39 377.93 l
	 317.41 383.40 l
	 313.76 383.16 l
cp p3
np
  317.39 377.93 m
	 321.08 377.93 l
	 321.06 383.40 l
	 317.41 383.40 l
cp p3
np
  321.08 377.93 m
	 324.78 377.75 l
	 324.71 383.16 l
	 321.06 383.40 l
cp p3
np
  324.78 377.75 m
	 328.46 377.38 l
	 328.36 382.70 l
	 324.71 383.16 l
cp p3
np
  328.46 377.38 m
	 332.15 376.87 l
	 332.00 382.03 l
	 328.36 382.70 l
cp p3
np
  332.15 376.87 m
	 335.82 376.22 l
	 335.62 381.18 l
	 332.00 382.03 l
cp p3
np
  335.82 376.22 m
	 339.49 375.47 l
	 339.24 380.18 l
	 335.62 381.18 l
cp p3
np
  339.49 375.47 m
	 343.14 374.66 l
	 342.84 379.10 l
	 339.24 380.18 l
cp p3
np
  343.14 374.66 m
	 346.79 373.81 l
	 346.43 377.99 l
	 342.84 379.10 l
cp p3
np
  346.79 373.81 m
	 350.43 372.95 l
	 350.01 376.88 l
	 346.43 377.99 l
cp p3
np
  350.43 372.95 m
	 354.06 372.10 l
	 353.59 375.80 l
	 350.01 376.88 l
cp p3
np
  251.94 366.45 m
	 255.54 366.87 l
	 256.48 369.51 l
	 252.94 369.02 l
cp p3
np
  255.54 366.87 m
	 259.14 367.35 l
	 260.03 370.05 l
	 256.48 369.51 l
cp p3
np
  259.14 367.35 m
	 262.74 367.87 l
	 263.57 370.66 l
	 260.03 370.05 l
cp p3
np
  262.74 367.87 m
	 266.35 368.45 l
	 267.12 371.34 l
	 263.57 370.66 l
cp p3
np
  248.33 366.06 m
	 251.94 366.45 l
	 252.94 369.02 l
	 249.40 368.58 l
cp p3
np
  365.59 366.65 m
	 369.26 366.08 l
	 368.52 369.08 l
	 364.91 369.76 l
cp p3
np
  369.26 366.08 m
	 372.92 365.55 l
	 372.13 368.45 l
	 368.52 369.08 l
cp p3
np
  372.92 365.55 m
	 376.59 365.06 l
	 375.73 367.87 l
	 372.13 368.45 l
cp p3
np
  361.91 367.25 m
	 365.59 366.65 l
	 364.91 369.76 l
	 361.30 370.49 l
cp p3
np
  380.25 364.61 m
	 383.91 364.20 l
	 382.94 366.87 l
	 379.34 367.35 l
cp p3
np
  383.91 364.20 m
	 387.58 363.82 l
	 386.54 366.45 l
	 382.94 366.87 l
cp p3
np
  387.58 363.82 m
	 391.24 363.48 l
	 390.14 366.06 l
	 386.54 366.45 l
cp p3
np
  376.59 365.06 m
	 380.25 364.61 l
	 379.34 367.35 l
	 375.73 367.87 l
cp p3
np
  347.17 369.90 m
	 350.86 369.22 l
	 350.43 372.95 l
	 346.79 373.81 l
cp p3
np
  350.86 369.22 m
	 354.55 368.55 l
	 354.06 372.10 l
	 350.43 372.95 l
cp p3
np
  354.55 368.55 m
	 358.23 367.89 l
	 357.68 371.27 l
	 354.06 372.10 l
cp p3
np
  358.23 367.89 m
	 361.91 367.25 l
	 361.30 370.49 l
	 357.68 371.27 l
cp p3
np
  261.89 365.06 m
	 265.55 365.55 l
	 266.35 368.45 l
	 262.74 367.87 l
cp p3
np
  265.55 365.55 m
	 269.22 366.08 l
	 269.95 369.08 l
	 266.35 368.45 l
cp p3
np
  269.22 366.08 m
	 272.89 366.65 l
	 273.56 369.76 l
	 269.95 369.08 l
cp p3
np
  272.89 366.65 m
	 276.56 367.25 l
	 277.18 370.49 l
	 273.56 369.76 l
cp p3
np
  276.56 367.25 m
	 280.24 367.89 l
	 280.80 371.27 l
	 277.18 370.49 l
cp p3
np
  280.24 367.89 m
	 283.92 368.55 l
	 284.42 372.10 l
	 280.80 371.27 l
cp p3
np
  283.92 368.55 m
	 287.61 369.22 l
	 288.05 372.95 l
	 284.42 372.10 l
cp p3
np
  287.61 369.22 m
	 291.31 369.90 l
	 291.69 373.81 l
	 288.05 372.95 l
cp p3
np
  291.31 369.90 m
	 295.01 370.56 l
	 295.33 374.66 l
	 291.69 373.81 l
cp p3
np
  295.01 370.56 m
	 298.72 371.18 l
	 298.99 375.47 l
	 295.33 374.66 l
cp p3
np
  298.72 371.18 m
	 302.44 371.75 l
	 302.66 376.22 l
	 298.99 375.47 l
cp p3
np
  302.44 371.75 m
	 306.16 372.24 l
	 306.33 376.87 l
	 302.66 376.22 l
cp p3
np
  306.16 372.24 m
	 309.89 372.63 l
	 310.01 377.38 l
	 306.33 376.87 l
cp p3
np
  309.89 372.63 m
	 313.63 372.90 l
	 313.70 377.75 l
	 310.01 377.38 l
cp p3
np
  313.63 372.90 m
	 317.37 373.03 l
	 317.39 377.93 l
	 313.70 377.75 l
cp p3
np
  317.37 373.03 m
	 321.11 373.03 l
	 321.08 377.93 l
	 317.39 377.93 l
cp p3
np
  321.11 373.03 m
	 324.85 372.90 l
	 324.78 377.75 l
	 321.08 377.93 l
cp p3
np
  324.85 372.90 m
	 328.58 372.63 l
	 328.46 377.38 l
	 324.78 377.75 l
cp p3
np
  328.58 372.63 m
	 332.31 372.24 l
	 332.15 376.87 l
	 328.46 377.38 l
cp p3
np
  332.31 372.24 m
	 336.04 371.75 l
	 335.82 376.22 l
	 332.15 376.87 l
cp p3
np
  336.04 371.75 m
	 339.75 371.18 l
	 339.49 375.47 l
	 335.82 376.22 l
cp p3
np
  339.75 371.18 m
	 343.46 370.56 l
	 343.14 374.66 l
	 339.49 375.47 l
cp p3
np
  343.46 370.56 m
	 347.17 369.90 l
	 346.79 373.81 l
	 343.14 374.66 l
cp p3
np
  247.24 363.48 m
	 250.90 363.82 l
	 251.94 366.45 l
	 248.33 366.06 l
cp p3
np
  250.90 363.82 m
	 254.56 364.20 l
	 255.54 366.87 l
	 251.94 366.45 l
cp p3
np
  254.56 364.20 m
	 258.22 364.61 l
	 259.14 367.35 l
	 255.54 366.87 l
cp p3
np
  258.22 364.61 m
	 261.89 365.06 l
	 262.74 367.87 l
	 259.14 367.35 l
cp p3
np
  358.81 364.58 m
	 362.55 364.06 l
	 361.91 367.25 l
	 358.23 367.89 l
cp p3
np
  362.55 364.06 m
	 366.29 363.56 l
	 365.59 366.65 l
	 361.91 367.25 l
cp p3
np
  366.29 363.56 m
	 370.02 363.08 l
	 369.26 366.08 l
	 365.59 366.65 l
cp p3
np
  370.02 363.08 m
	 373.75 362.64 l
	 372.92 365.55 l
	 369.26 366.08 l
cp p3
np
  373.75 362.64 m
	 377.48 362.22 l
	 376.59 365.06 l
	 372.92 365.55 l
cp p3
np
  377.48 362.22 m
	 381.20 361.83 l
	 380.25 364.61 l
	 376.59 365.06 l
cp p3
np
  381.20 361.83 m
	 384.93 361.48 l
	 383.91 364.20 l
	 380.25 364.61 l
cp p3
np
  384.93 361.48 m
	 388.65 361.15 l
	 387.58 363.82 l
	 383.91 364.20 l
cp p3
np
  388.65 361.15 m
	 392.37 360.85 l
	 391.24 363.48 l
	 387.58 363.82 l
cp p3
np
  343.81 366.71 m
	 347.57 366.19 l
	 347.17 369.90 l
	 343.46 370.56 l
cp p3
np
  347.57 366.19 m
	 351.32 365.66 l
	 350.86 369.22 l
	 347.17 369.90 l
cp p3
np
  351.32 365.66 m
	 355.07 365.12 l
	 354.55 368.55 l
	 350.86 369.22 l
cp p3
np
  355.07 365.12 m
	 358.81 364.58 l
	 358.23 367.89 l
	 354.55 368.55 l
cp p3
np
  249.83 361.15 m
	 253.55 361.48 l
	 254.56 364.20 l
	 250.90 363.82 l
cp p3
np
  253.55 361.48 m
	 257.27 361.83 l
	 258.22 364.61 l
	 254.56 364.20 l
cp p3
np
  257.27 361.83 m
	 261.00 362.22 l
	 261.89 365.06 l
	 258.22 364.61 l
cp p3
np
  261.00 362.22 m
	 264.73 362.64 l
	 265.55 365.55 l
	 261.89 365.06 l
cp p3
np
  264.73 362.64 m
	 268.46 363.08 l
	 269.22 366.08 l
	 265.55 365.55 l
cp p3
np
  268.46 363.08 m
	 272.19 363.56 l
	 272.89 366.65 l
	 269.22 366.08 l
cp p3
np
  272.19 363.56 m
	 275.92 364.06 l
	 276.56 367.25 l
	 272.89 366.65 l
cp p3
np
  275.92 364.06 m
	 279.66 364.58 l
	 280.24 367.89 l
	 276.56 367.25 l
cp p3
np
  279.66 364.58 m
	 283.41 365.12 l
	 283.92 368.55 l
	 280.24 367.89 l
cp p3
np
  283.41 365.12 m
	 287.15 365.66 l
	 287.61 369.22 l
	 283.92 368.55 l
cp p3
np
  287.15 365.66 m
	 290.91 366.19 l
	 291.31 369.90 l
	 287.61 369.22 l
cp p3
np
  290.91 366.19 m
	 294.67 366.71 l
	 295.01 370.56 l
	 291.31 369.90 l
cp p3
np
  294.67 366.71 m
	 298.44 367.19 l
	 298.72 371.18 l
	 295.01 370.56 l
cp p3
np
  298.44 367.19 m
	 302.21 367.63 l
	 302.44 371.75 l
	 298.72 371.18 l
cp p3
np
  302.21 367.63 m
	 305.99 368.01 l
	 306.16 372.24 l
	 302.44 371.75 l
cp p3
np
  305.99 368.01 m
	 309.77 368.30 l
	 309.89 372.63 l
	 306.16 372.24 l
cp p3
np
  309.77 368.30 m
	 313.55 368.50 l
	 313.63 372.90 l
	 309.89 372.63 l
cp p3
np
  313.55 368.50 m
	 317.34 368.61 l
	 317.37 373.03 l
	 313.63 372.90 l
cp p3
np
  317.34 368.61 m
	 321.13 368.61 l
	 321.11 373.03 l
	 317.37 373.03 l
cp p3
np
  321.13 368.61 m
	 324.92 368.50 l
	 324.85 372.90 l
	 321.11 373.03 l
cp p3
np
  324.92 368.50 m
	 328.71 368.30 l
	 328.58 372.63 l
	 324.85 372.90 l
cp p3
np
  328.71 368.30 m
	 332.49 368.01 l
	 332.31 372.24 l
	 328.58 372.63 l
cp p3
np
  332.49 368.01 m
	 336.27 367.63 l
	 336.04 371.75 l
	 332.31 372.24 l
cp p3
np
  336.27 367.63 m
	 340.04 367.19 l
	 339.75 371.18 l
	 336.04 371.75 l
cp p3
np
  340.04 367.19 m
	 343.81 366.71 l
	 343.46 370.56 l
	 339.75 371.18 l
cp p3
np
  246.10 360.85 m
	 249.83 361.15 l
	 250.90 363.82 l
	 247.24 363.48 l
cp p3
np
  340.34 363.42 m
	 344.17 363.04 l
	 343.81 366.71 l
	 340.04 367.19 l
cp p3
np
  347.99 362.63 m
	 351.80 362.20 l
	 351.32 365.66 l
	 347.57 366.19 l
cp p3
np
  351.80 362.20 m
	 355.61 361.76 l
	 355.07 365.12 l
	 351.32 365.66 l
cp p3
np
  355.61 361.76 m
	 359.42 361.32 l
	 358.81 364.58 l
	 355.07 365.12 l
cp p3
np
  359.42 361.32 m
	 363.22 360.89 l
	 362.55 364.06 l
	 358.81 364.58 l
cp p3
np
  363.22 360.89 m
	 367.02 360.48 l
	 366.29 363.56 l
	 362.55 364.06 l
cp p3
np
  367.02 360.48 m
	 370.81 360.08 l
	 370.02 363.08 l
	 366.29 363.56 l
cp p3
np
  370.81 360.08 m
	 374.61 359.70 l
	 373.75 362.64 l
	 370.02 363.08 l
cp p3
np
  374.61 359.70 m
	 378.40 359.34 l
	 377.48 362.22 l
	 373.75 362.64 l
cp p3
np
  378.40 359.34 m
	 382.18 359.01 l
	 381.20 361.83 l
	 377.48 362.22 l
cp p3
np
  382.18 359.01 m
	 385.97 358.70 l
	 384.93 361.48 l
	 381.20 361.83 l
cp p3
np
  385.97 358.70 m
	 389.76 358.41 l
	 388.65 361.15 l
	 384.93 361.48 l
cp p3
np
  389.76 358.41 m
	 393.54 358.15 l
	 392.37 360.85 l
	 388.65 361.15 l
cp p3
np
  344.17 363.04 m
	 347.99 362.63 l
	 347.57 366.19 l
	 343.81 366.71 l
cp p3
np
  244.93 358.15 m
	 248.72 358.41 l
	 249.83 361.15 l
	 246.10 360.85 l
cp p3
np
  248.72 358.41 m
	 252.50 358.70 l
	 253.55 361.48 l
	 249.83 361.15 l
cp p3
np
  252.50 358.70 m
	 256.29 359.01 l
	 257.27 361.83 l
	 253.55 361.48 l
cp p3
np
  256.29 359.01 m
	 260.08 359.34 l
	 261.00 362.22 l
	 257.27 361.83 l
cp p3
np
  260.08 359.34 m
	 263.87 359.70 l
	 264.73 362.64 l
	 261.00 362.22 l
cp p3
np
  263.87 359.70 m
	 267.66 360.08 l
	 268.46 363.08 l
	 264.73 362.64 l
cp p3
np
  267.66 360.08 m
	 271.46 360.48 l
	 272.19 363.56 l
	 268.46 363.08 l
cp p3
np
  271.46 360.48 m
	 275.26 360.89 l
	 275.92 364.06 l
	 272.19 363.56 l
cp p3
np
  275.26 360.89 m
	 279.06 361.32 l
	 279.66 364.58 l
	 275.92 364.06 l
cp p3
np
  279.06 361.32 m
	 282.86 361.76 l
	 283.41 365.12 l
	 279.66 364.58 l
cp p3
np
  282.86 361.76 m
	 286.67 362.20 l
	 287.15 365.66 l
	 283.41 365.12 l
cp p3
np
  286.67 362.20 m
	 290.49 362.63 l
	 290.91 366.19 l
	 287.15 365.66 l
cp p3
np
  290.49 362.63 m
	 294.31 363.04 l
	 294.67 366.71 l
	 290.91 366.19 l
cp p3
np
  294.31 363.04 m
	 298.13 363.42 l
	 298.44 367.19 l
	 294.67 366.71 l
cp p3
np
  298.13 363.42 m
	 301.96 363.76 l
	 302.21 367.63 l
	 298.44 367.19 l
cp p3
np
  301.96 363.76 m
	 305.80 364.05 l
	 305.99 368.01 l
	 302.21 367.63 l
cp p3
np
  305.80 364.05 m
	 309.63 364.28 l
	 309.77 368.30 l
	 305.99 368.01 l
cp p3
np
  309.63 364.28 m
	 313.47 364.43 l
	 313.55 368.50 l
	 309.77 368.30 l
cp p3
np
  313.47 364.43 m
	 317.32 364.51 l
	 317.34 368.61 l
	 313.55 368.50 l
cp p3
np
  317.32 364.51 m
	 321.16 364.51 l
	 321.13 368.61 l
	 317.34 368.61 l
cp p3
np
  321.16 364.51 m
	 325.00 364.43 l
	 324.92 368.50 l
	 321.13 368.61 l
cp p3
np
  325.00 364.43 m
	 328.84 364.28 l
	 328.71 368.30 l
	 324.92 368.50 l
cp p3
np
  328.84 364.28 m
	 332.68 364.05 l
	 332.49 368.01 l
	 328.71 368.30 l
cp p3
np
  332.68 364.05 m
	 336.51 363.76 l
	 336.27 367.63 l
	 332.49 368.01 l
cp p3
np
  336.51 363.76 m
	 340.34 363.42 l
	 340.04 367.19 l
	 336.27 367.63 l
cp p3
ep
%%Trailer
%%Pages: 1
%%EOF
