%!PS-Adobe-3.0
%%DocumentNeededResources: font Helvetica
%%+ font Helvetica-Bold
%%+ font Helvetica-Oblique
%%+ font Helvetica-BoldOblique
%%+ font Symbol
%%DocumentMedia: a4 595 841 0 () ()
%%Title: R Graphics Output
%%Creator: R Software
%%Pages: (atend)
%%Orientation: Landscape
%%BoundingBox: 18 18 577 824
%%EndComments
%%BeginProlog
/bp  { gs 595.00 0 translate 90 rotate gs } def
% begin .ps.prolog
/gs  { gsave } def
/gr  { grestore } def
/ep  { showpage gr gr } def
/m   { moveto } def
/l   { lineto } def
/np  { newpath } def
/cp  { closepath } def
/f   { fill } def
/o   { stroke } def
/c   { newpath 0 360 arc } def
/r   { 3 index 3 index moveto 1 index 4 -1 roll
       lineto exch 1 index lineto lineto closepath } def
/p1  { stroke } def
/p2  { gsave bg setrgbcolor fill grestore newpath } def
/p3  { gsave bg setrgbcolor fill grestore stroke } def
/t   { 6 -2 roll moveto gsave rotate
       ps mul neg 0 2 1 roll rmoveto
       1 index stringwidth pop
       mul neg 0 rmoveto show grestore } def
/cl  { grestore gsave newpath 3 index 3 index moveto 1 index
       4 -1 roll lineto  exch 1 index lineto lineto
       closepath clip newpath } def
/rgb { setrgbcolor } def
/s   { scalefont setfont } def
/R   { /Font1 findfont } def
/B   { /Font2 findfont } def
/I   { /Font3 findfont } def
/BI  { /Font4 findfont } def
/S   { /Font5 findfont } def
1 setlinecap 1 setlinejoin
% end   .ps.prolog
%%IncludeResource: font Helvetica
/Helvetica findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font1 exch definefont pop
%%IncludeResource: font Helvetica-Bold
/Helvetica-Bold findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font2 exch definefont pop
%%IncludeResource: font Helvetica-Oblique
/Helvetica-Oblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font3 exch definefont pop
%%IncludeResource: font Helvetica-BoldOblique
/Helvetica-BoldOblique findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font4 exch definefont pop
%%IncludeResource: font Symbol
/Symbol findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  currentdict
  end
/Font5 exch definefont pop
%%EndProlog
%%Page: 1 1
bp
18.00 18.00 823.89 577.28 cl
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
238.15 91.44 m
633.33 91.44 l
o
np
238.15 91.44 m
238.15 84.24 l
o
np
317.19 91.44 m
317.19 84.24 l
o
np
396.22 91.44 m
396.22 84.24 l
o
np
475.26 91.44 m
475.26 84.24 l
o
np
554.29 91.44 m
554.29 84.24 l
o
np
633.33 91.44 m
633.33 84.24 l
o
/ps 12 def R 12 s
238.15 65.52 (540000) 0.50 0.00 0.00 t
317.19 65.52 (540200) 0.50 0.00 0.00 t
396.22 65.52 (540400) 0.50 0.00 0.00 t
475.26 65.52 (540600) 0.50 0.00 0.00 t
554.29 65.52 (540800) 0.50 0.00 0.00 t
633.33 65.52 (541000) 0.50 0.00 0.00 t
np
221.95 107.25 m
221.95 502.43 l
o
np
221.95 107.25 m
214.75 107.25 l
o
np
221.95 186.28 m
214.75 186.28 l
o
np
221.95 265.32 m
214.75 265.32 l
o
np
221.95 344.36 m
214.75 344.36 l
o
np
221.95 423.39 m
214.75 423.39 l
o
np
221.95 502.43 m
214.75 502.43 l
o
204.67 107.25 (1794000) 0.50 0.00 90.00 t
204.67 186.28 (1794200) 0.50 0.00 90.00 t
204.67 265.32 (1794400) 0.50 0.00 90.00 t
204.67 344.36 (1794600) 0.50 0.00 90.00 t
204.67 423.39 (1794800) 0.50 0.00 90.00 t
204.67 502.43 (1795000) 0.50 0.00 90.00 t
np
221.95 91.44 m
648.74 91.44 l
648.74 518.24 l
221.95 518.24 l
221.95 91.44 l
o
221.95 91.44 648.74 518.24 cl
/bg { 1.0000 0.0000 0.0000 } def
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
  283.99 502.43 m
	 341.29 502.43 l
	 346.43 470.81 l
	 293.08 462.91 l
cp p3
/bg { 1.0000 0.0902 0.0000 } def
np
  387.53 502.43 m
	 422.70 502.43 l
	 417.17 443.15 l
	 385.55 443.15 l
	 385.95 458.96 l
cp p3
/bg { 1.0000 0.1804 0.0000 } def
np
  345.64 458.96 m
	 346.43 443.15 l
	 348.01 423.39 l
	 299.80 431.30 l
	 297.82 439.20 l
	 335.76 451.05 l
cp p3
/bg { 1.0000 0.2745 0.0000 } def
np
  341.29 502.43 m
	 387.53 502.43 l
	 385.95 458.96 l
	 381.21 458.96 l
	 363.82 458.96 l
	 362.63 490.57 l
	 357.10 490.57 l
	 358.28 466.86 l
	 361.05 455.01 l
	 380.81 455.01 l
	 379.23 419.44 l
	 370.93 419.44 l
	 365.79 447.10 l
	 346.43 443.15 l
	 345.64 458.96 l
	 346.03 470.81 l
cp p3
/bg { 1.0000 0.3647 0.0000 } def
np
  385.55 443.15 m
	 417.17 443.15 l
	 414.01 407.58 l
	 395.43 407.58 l
	 383.18 415.49 l
cp p3
/bg { 1.0000 0.4549 0.0000 } def
np
  422.70 502.43 m
	 457.87 502.43 l
	 457.08 403.63 l
	 414.01 407.58 l
	 417.17 443.15 l
cp p3
/bg { 1.0000 0.5451 0.0000 } def
np
  457.87 502.43 m
	 496.20 502.43 l
	 500.55 439.20 l
	 509.24 439.20 l
	 513.20 399.68 l
	 457.08 403.63 l
	 457.48 451.05 l
cp p3
/bg { 1.0000 0.6353 0.0000 } def
np
  299.80 427.34 m
	 301.38 431.30 l
	 329.04 427.34 l
	 335.76 395.73 l
	 306.12 395.73 l
cp p3
/bg { 1.0000 0.7255 0.0000 } def
np
  306.12 395.73 m
	 335.76 395.73 l
	 336.55 379.92 l
	 309.68 379.92 l
cp p3
/bg { 1.0000 0.8196 0.0000 } def
np
  309.68 379.92 m
	 319.56 379.92 l
	 329.44 332.50 l
	 321.93 328.55 l
	 321.93 332.50 l
	 322.32 336.45 l
	 323.11 344.36 l
	 323.11 348.31 l
	 322.32 352.26 l
	 319.16 356.21 l
	 314.42 356.21 l
cp p3
/bg { 1.0000 0.9098 0.0000 } def
np
  401.36 292.98 m
	 398.20 344.36 l
	 456.68 348.31 l
	 456.29 296.93 l
cp p3
/bg { 1.0000 1.0000 0.0000 } def
np
  389.50 403.63 m
	 456.68 399.68 l
	 456.68 348.31 l
	 398.20 344.36 l
cp p3
/bg { 0.9098 1.0000 0.0000 } def
np
  359.07 348.31 m
	 398.20 344.36 l
	 401.36 292.98 l
	 385.55 289.03 l
cp p3
/bg { 0.8196 1.0000 0.0000 } def
np
  329.04 427.34 m
	 373.70 419.44 l
	 374.09 419.44 l
	 389.50 403.63 l
	 398.20 344.36 l
	 359.07 348.31 l
	 355.91 352.26 l
	 342.87 379.92 l
	 336.55 379.92 l
	 335.76 395.73 l
cp p3
/bg { 0.7255 1.0000 0.0000 } def
np
  322.72 328.55 m
	 329.04 328.55 l
	 340.50 281.13 l
	 331.41 281.13 l
	 330.62 285.08 l
	 328.25 285.08 l
cp p3
/bg { 0.6353 1.0000 0.0000 } def
np
  332.20 277.18 m
	 344.06 277.18 l
	 357.10 281.13 l
	 357.89 273.22 l
	 387.13 281.13 l
	 411.24 202.09 l
	 350.38 186.28 l
	 332.20 273.22 l
cp p3
/bg { 0.5451 1.0000 0.0000 } def
np
  388.71 285.08 m
	 419.54 289.03 l
	 450.36 292.98 l
	 478.42 296.93 l
	 486.72 221.85 l
	 482.37 221.85 l
	 422.30 202.09 l
	 420.72 206.04 l
	 416.38 206.04 l
cp p3
/bg { 0.4549 1.0000 0.0000 } def
np
  427.84 107.25 m
	 427.84 123.05 l
	 429.02 142.81 l
	 430.60 154.67 l
	 432.58 170.48 l
	 430.21 186.28 l
	 425.07 198.14 l
	 422.30 202.09 l
	 474.86 217.90 l
	 488.69 217.90 l
	 491.07 198.14 l
	 492.25 194.19 l
	 535.72 186.28 l
	 530.98 166.52 l
	 528.21 127.01 l
	 527.82 107.25 l
cp p3
/bg { 0.3647 1.0000 0.0000 } def
np
  238.54 466.86 m
	 238.15 502.43 l
	 278.46 502.43 l
	 285.18 466.86 l
cp p3
/bg { 0.2745 1.0000 0.0000 } def
np
  238.94 372.02 m
	 238.15 466.86 l
	 265.42 466.86 l
	 282.80 379.92 l
	 273.72 375.97 l
	 255.14 375.97 l
cp p3
/bg { 0.1804 1.0000 0.0000 } def
np
  265.42 466.86 m
	 278.85 466.86 l
	 296.24 379.92 l
	 282.80 379.92 l
cp p3
/bg { 0.0902 1.0000 0.0000 } def
np
  296.24 379.92 m
	 278.85 466.86 l
	 286.76 466.86 l
	 296.24 423.39 l
	 301.77 379.92 l
cp p3
/bg { 0.0000 1.0000 0.0000 } def
np
  238.54 340.40 m
	 263.44 344.36 l
	 275.30 257.42 l
	 238.54 253.46 l
cp p3
/bg { 0.0000 1.0000 0.0902 } def
np
  271.74 285.08 m
	 307.70 292.98 l
	 327.46 261.37 l
	 275.30 257.42 l
cp p3
/bg { 0.0000 1.0000 0.1804 } def
np
  238.54 253.46 m
	 275.30 257.42 l
	 278.06 229.75 l
	 238.54 225.80 l
cp p3
/bg { 0.0000 1.0000 0.2745 } def
np
  275.30 257.42 m
	 327.46 261.37 l
	 334.57 233.71 l
	 278.06 229.75 l
cp p3
/bg { 0.0000 1.0000 0.3647 } def
np
  238.54 225.80 m
	 278.06 229.75 l
	 282.80 198.14 l
	 238.15 190.24 l
cp p3
/bg { 0.0000 1.0000 0.4549 } def
np
  278.06 229.75 m
	 334.57 233.71 l
	 344.45 190.24 l
	 319.56 186.28 l
	 317.98 194.19 l
	 313.23 198.14 l
	 304.94 202.09 l
	 301.77 209.99 l
	 281.22 206.04 l
cp p3
/bg { 0.0000 1.0000 0.5451 } def
np
  318.37 182.33 m
	 345.24 186.28 l
	 351.57 158.62 l
	 316.79 158.62 l
	 314.42 174.43 l
cp p3
/bg { 0.0000 1.0000 0.6353 } def
np
  238.15 190.24 m
	 273.72 194.19 l
	 274.11 182.33 l
	 280.83 178.38 l
	 283.20 182.33 l
	 283.20 174.43 l
	 238.15 174.43 l
cp p3
/bg { 0.0000 1.0000 0.7255 } def
np
  238.15 174.43 m
	 283.20 174.43 l
	 286.76 154.67 l
	 237.75 150.72 l
cp p3
/bg { 0.0000 1.0000 0.8196 } def
np
  237.75 150.72 m
	 286.76 154.67 l
	 293.87 107.25 l
	 238.54 107.25 l
cp p3
/bg { 0.0000 1.0000 0.9098 } def
np
  293.87 107.25 m
	 286.76 154.67 l
	 287.94 154.67 l
	 316.79 158.62 l
	 351.57 158.62 l
	 361.45 107.25 l
cp p3
/bg { 0.0000 1.0000 1.0000 } def
np
  350.38 186.28 m
	 360.26 186.28 l
	 364.61 158.62 l
	 365.00 150.72 l
	 357.89 150.72 l
cp p3
/bg { 0.0000 0.9098 1.0000 } def
np
  360.26 186.28 m
	 411.24 202.09 l
	 412.82 202.09 l
	 423.09 186.28 l
	 426.26 174.43 l
	 425.47 154.67 l
	 367.77 146.77 l
	 365.00 150.72 l
	 364.61 158.62 l
cp p3
/bg { 0.0000 0.8196 1.0000 } def
np
  375.28 107.25 m
	 367.77 146.77 l
	 425.47 154.67 l
	 423.49 134.91 l
	 421.12 127.01 l
	 419.93 107.25 l
cp p3
/bg { 0.0000 0.7255 1.0000 } def
np
  367.37 107.25 m
	 363.03 123.05 l
	 359.87 142.81 l
	 363.03 146.77 l
	 367.77 130.96 l
	 372.91 107.25 l
cp p3
/bg { 0.0000 0.6353 1.0000 } def
np
  478.42 296.93 m
	 503.71 296.93 l
	 510.43 249.51 l
	 487.51 245.56 l
	 491.07 225.80 l
	 486.72 221.85 l
cp p3
/bg { 0.0000 0.5451 1.0000 } def
np
  503.71 296.93 m
	 519.12 300.89 l
	 526.63 249.51 l
	 510.43 249.51 l
cp p3
/bg { 0.0000 0.4549 1.0000 } def
np
  519.12 300.89 m
	 550.74 300.89 l
	 561.01 300.89 l
	 570.10 300.89 l
	 560.22 285.08 l
	 562.59 277.18 l
	 577.61 273.22 l
	 563.78 253.46 l
	 526.63 249.51 l
cp p3
/bg { 0.0000 0.3647 1.0000 } def
np
  591.84 292.98 m
	 608.04 292.98 l
	 616.34 289.03 l
	 624.64 292.98 l
	 624.64 253.46 l
	 569.71 249.51 l
cp p3
/bg { 0.0000 0.2745 1.0000 } def
np
  569.71 249.51 m
	 624.64 253.46 l
	 626.22 209.99 l
	 548.37 213.95 l
	 558.25 229.75 l
cp p3
/bg { 0.0000 0.1804 1.0000 } def
np
  548.37 213.95 m
	 626.22 209.99 l
	 626.61 150.72 l
	 547.18 154.67 l
	 547.18 198.14 l
	 543.62 202.09 l
cp p3
/bg { 0.0000 0.0902 1.0000 } def
np
  555.48 107.25 m
	 555.88 127.01 l
	 560.22 138.86 l
	 563.78 154.67 l
	 626.61 150.72 l
	 625.82 134.91 l
	 626.61 107.25 l
cp p3
/bg { 0.0000 0.0000 1.0000 } def
np
  488.69 217.90 m
	 493.83 221.85 l
	 496.60 213.95 l
	 501.74 209.99 l
	 502.92 198.14 l
	 491.07 198.14 l
cp p3
/bg { 0.0902 0.0000 1.0000 } def
np
  501.74 209.99 m
	 522.68 206.04 l
	 528.61 209.99 l
	 534.93 225.80 l
	 551.92 229.75 l
	 543.62 209.99 l
	 535.33 190.24 l
	 502.92 198.14 l
cp p3
/bg { 0.1804 0.0000 1.0000 } def
np
  528.61 249.51 m
	 563.78 253.46 l
	 557.85 233.71 l
	 549.55 233.71 l
	 548.76 237.66 l
	 538.49 237.66 l
	 538.09 245.56 l
	 530.19 245.56 l
cp p3
/bg { 0.2745 0.0000 1.0000 } def
np
  459.06 399.68 m
	 463.01 403.63 l
	 465.38 403.63 l
	 486.72 399.68 l
	 486.32 395.73 l
	 487.51 375.97 l
	 459.45 372.02 l
cp p3
/bg { 0.3647 0.0000 1.0000 } def
np
  459.45 372.02 m
	 487.51 375.97 l
	 486.72 348.31 l
	 459.85 348.31 l
cp p3
/bg { 0.4549 0.0000 1.0000 } def
np
  486.72 399.68 m
	 511.22 399.68 l
	 511.22 304.84 l
	 486.72 300.89 l
	 486.72 348.31 l
	 487.51 375.97 l
	 486.32 395.73 l
cp p3
/bg { 0.5451 0.0000 1.0000 } def
np
  511.22 399.68 m
	 521.89 395.73 l
	 521.49 383.87 l
	 529.79 383.87 l
	 528.61 304.84 l
	 511.22 304.84 l
cp p3
/bg { 0.6353 0.0000 1.0000 } def
np
  528.61 304.84 m
	 529.40 348.31 l
	 555.48 348.31 l
	 555.48 312.74 l
	 547.18 312.74 l
	 546.39 308.79 l
	 535.33 308.79 l
	 532.56 304.84 l
cp p3
/bg { 0.7255 0.0000 1.0000 } def
np
  557.06 395.73 m
	 597.76 395.73 l
	 598.95 352.26 l
	 555.88 348.31 l
	 555.48 383.87 l
cp p3
/bg { 0.8196 0.0000 1.0000 } def
np
  555.88 348.31 m
	 598.95 352.26 l
	 604.48 320.65 l
	 588.28 320.65 l
	 587.09 308.79 l
	 559.43 308.79 l
	 555.48 312.74 l
	 555.48 348.31 l
cp p3
/bg { 0.9098 0.0000 1.0000 } def
np
  616.73 308.79 m
	 611.60 324.60 l
	 609.22 352.26 l
	 608.04 375.97 l
	 604.48 379.92 l
	 604.09 391.78 l
	 624.64 391.78 l
	 624.64 312.74 l
cp p3
/bg { 1.0000 0.0000 1.0000 } def
np
  496.20 502.43 m
	 518.73 502.43 l
	 521.49 439.20 l
	 500.15 439.20 l
cp p3
/bg { 1.0000 0.0000 0.9098 } def
np
  513.20 439.20 m
	 521.49 439.20 l
	 519.52 486.62 l
	 535.72 482.67 l
	 547.18 399.68 l
	 516.75 403.63 l
cp p3
/bg { 1.0000 0.0000 0.8196 } def
np
  518.73 502.43 m
	 539.28 502.43 l
	 540.46 494.52 l
	 540.86 486.62 l
	 549.55 486.62 l
	 556.67 466.86 l
	 538.49 462.91 l
	 535.72 482.67 l
	 519.52 486.62 l
cp p3
/bg { 1.0000 0.0000 0.7255 } def
np
  539.28 502.43 m
	 601.72 502.43 l
	 604.48 470.81 l
	 556.67 466.86 l
	 549.55 486.62 l
	 540.86 486.62 l
	 540.46 494.52 l
cp p3
/bg { 1.0000 0.0000 0.6353 } def
np
  604.48 470.81 m
	 604.48 435.25 l
	 600.93 435.25 l
	 548.37 427.34 l
	 544.81 466.86 l
	 556.67 466.86 l
cp p3
/bg { 1.0000 0.0000 0.5451 } def
np
  548.37 427.34 m
	 576.82 431.30 l
	 600.93 435.25 l
	 604.48 435.25 l
	 600.14 395.73 l
	 548.76 399.68 l
cp p3
/bg { 1.0000 0.0000 0.4549 } def
np
  604.09 502.43 m
	 625.03 502.43 l
	 625.03 474.77 l
	 607.64 474.77 l
cp p3
/bg { 1.0000 0.0000 0.3647 } def
np
  607.64 474.77 m
	 625.03 474.77 l
	 625.03 415.49 l
	 604.48 415.49 l
	 604.48 435.25 l
cp p3
/bg { 1.0000 0.0000 0.2745 } def
np
  604.48 415.49 m
	 625.03 415.49 l
	 624.64 391.78 l
	 604.09 391.78 l
	 601.32 403.63 l
cp p3
/bg { 1.0000 0.0000 0.1804 } def
np
  543.23 202.09 m
	 545.21 198.14 l
	 547.18 198.14 l
	 547.18 154.67 l
	 533.35 154.67 l
	 535.72 178.38 l
cp p3
/bg { 1.0000 0.0000 0.0902 } def
np
  293.08 462.91 m
	 346.43 470.81 l
	 345.64 458.96 l
	 335.76 451.05 l
	 297.82 439.20 l
	 295.85 451.05 l
cp p3
/ps 12 def R 12 s
316.20 480.43 (1) 0.50 0.00 0.00 t
399.78 465.81 (2) 0.50 0.00 0.00 t
328.91 437.07 (3) 0.50 0.00 0.00 t
364.61 458.20 (4) 0.50 0.00 0.00 t
399.07 419.38 (5) 0.50 0.00 0.00 t
433.76 447.74 (6) 0.50 0.00 0.00 t
484.52 444.10 (7) 0.50 0.00 0.00 t
314.42 411.38 (8) 0.50 0.00 0.00 t
322.03 383.72 (9) 0.50 0.00 0.00 t
320.63 345.64 (10) 0.50 0.00 0.00 t
428.13 316.43 (11) 0.50 0.00 0.00 t
425.27 369.78 (12) 0.50 0.00 0.00 t
386.05 314.57 (13) 0.50 0.00 0.00 t
359.47 382.82 (14) 0.50 0.00 0.00 t
330.42 294.15 (15) 0.50 0.00 0.00 t
359.03 252.32 (16) 0.50 0.00 0.00 t
440.61 242.66 (17) 0.50 0.00 0.00 t
468.44 164.64 (18) 0.50 0.00 0.00 t
260.08 480.54 (19) 0.50 0.00 0.00 t
259.03 402.16 (20) 0.50 0.00 0.00 t
280.83 419.17 (21) 0.50 0.00 0.00 t
291.97 419.17 (22) 0.50 0.00 0.00 t
253.96 294.81 (23) 0.50 0.00 0.00 t
295.55 269.99 (24) 0.50 0.00 0.00 t
257.61 237.50 (25) 0.50 0.00 0.00 t
303.85 241.46 (26) 0.50 0.00 0.00 t
259.39 206.76 (27) 0.50 0.00 0.00 t
310.64 201.50 (28) 0.50 0.00 0.00 t
329.28 167.95 (29) 0.50 0.00 0.00 t
267.34 178.23 (30) 0.50 0.00 0.00 t
261.47 159.46 (31) 0.50 0.00 0.00 t
264.23 125.87 (32) 0.50 0.00 0.00 t
316.40 136.08 (33) 0.50 0.00 0.00 t
359.63 162.42 (34) 0.50 0.00 0.00 t
395.17 169.45 (35) 0.50 0.00 0.00 t
405.51 125.54 (36) 0.50 0.00 0.00 t
365.66 122.24 (37) 0.50 0.00 0.00 t
492.98 251.99 (38) 0.50 0.00 0.00 t
514.97 270.11 (39) 0.50 0.00 0.00 t
554.65 278.34 (40) 0.50 0.00 0.00 t
605.87 274.27 (41) 0.50 0.00 0.00 t
585.43 227.12 (42) 0.50 0.00 0.00 t
573.20 184.16 (43) 0.50 0.00 0.00 t
587.77 127.30 (44) 0.50 0.00 0.00 t
495.81 205.89 (45) 0.50 0.00 0.00 t
527.72 205.89 (46) 0.50 0.00 0.00 t
544.41 237.88 (47) 0.50 0.00 0.00 t
472.49 388.80 (48) 0.50 0.00 0.00 t
473.38 357.05 (49) 0.50 0.00 0.00 t
493.78 356.62 (50) 0.50 0.00 0.00 t
520.70 358.04 (51) 0.50 0.00 0.00 t
541.30 314.57 (52) 0.50 0.00 0.00 t
573.03 371.08 (53) 0.50 0.00 0.00 t
575.63 323.46 (54) 0.50 0.00 0.00 t
612.93 350.72 (55) 0.50 0.00 0.00 t
509.14 466.71 (56) 0.50 0.00 0.00 t
525.64 437.82 (57) 0.50 0.00 0.00 t
537.70 481.64 (58) 0.50 0.00 0.00 t
561.86 483.08 (59) 0.50 0.00 0.00 t
576.62 446.29 (60) 0.50 0.00 0.00 t
579.92 416.65 (61) 0.50 0.00 0.00 t
615.45 484.49 (62) 0.50 0.00 0.00 t
613.33 439.05 (63) 0.50 0.00 0.00 t
611.91 399.53 (64) 0.50 0.00 0.00 t
541.98 176.91 (65) 0.50 0.00 0.00 t
319.10 451.56 (66) 0.50 0.00 0.00 t
ep
%%Trailer
%%Pages: 1
%%EOF
