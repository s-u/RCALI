%!PS-Adobe-3.0 EPSF-3.0
%%DocumentNeededResources: font Times-Roman
%%+ font Times-Bold
%%+ font Times-Italic
%%+ font Times-BoldItalic
%%+ font Symbol
%%Title: R Graphics Output
%%Creator: R Software
%%Pages: (atend)
%%BoundingBox: 118 277 478 565
%%EndComments
%%BeginProlog
/bp  { gs gs } def
% begin .ps.prolog
/gs  { gsave } def
/gr  { grestore } def
/ep  { showpage gr gr } def
/m   { moveto } def
/l   { lineto } def
/np  { newpath } def
/cp  { closepath } def
/f   { fill } def
/o   { stroke } def
/c   { newpath 0 360 arc } def
/r   { 3 index 3 index moveto 1 index 4 -1 roll
       lineto exch 1 index lineto lineto closepath } def
/p1  { stroke } def
/p2  { gsave bg setrgbcolor fill grestore newpath } def
/p3  { gsave bg setrgbcolor fill grestore stroke } def
/t   { 6 -2 roll moveto gsave rotate
       ps mul neg 0 2 1 roll rmoveto
       1 index stringwidth pop
       mul neg 0 rmoveto show grestore } def
/cl  { grestore gsave newpath 3 index 3 index moveto 1 index
       4 -1 roll lineto  exch 1 index lineto lineto
       closepath clip newpath } def
/rgb { setrgbcolor } def
/s   { scalefont setfont } def
/R   { /Font1 findfont } def
/B   { /Font2 findfont } def
/I   { /Font3 findfont } def
/BI  { /Font4 findfont } def
/S   { /Font5 findfont } def
1 setlinecap 1 setlinejoin
% end   .ps.prolog
%%IncludeResource: font Times-Roman
/Times-Roman findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font1 exch definefont pop
%%IncludeResource: font Times-Bold
/Times-Bold findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font2 exch definefont pop
%%IncludeResource: font Times-Italic
/Times-Italic findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font3 exch definefont pop
%%IncludeResource: font Times-BoldItalic
/Times-BoldItalic findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  /Encoding ISOLatin1Encoding def
  currentdict
  end
/Font4 exch definefont pop
%%IncludeResource: font Symbol
/Symbol findfont
dup length dict begin
  {1 index /FID ne {def} {pop pop} ifelse} forall
  currentdict
  end
/Font5 exch definefont pop
%%EndProlog
%%Page: 1 1
bp
171.76 344.26 463.12 550.42 cl
/ps 11 def R 11 s
0.0000 0.0000 0.0000 rgb
182.55 460.89 (1) 0.50 0.00 0.00 t
249.99 440.78 (1) 0.50 0.00 0.00 t
281.35 435.69 (1) 0.50 0.00 0.00 t
302.01 419.52 (1) 0.50 0.00 0.00 t
317.44 417.42 (1) 0.50 0.00 0.00 t
329.76 414.37 (1) 0.50 0.00 0.00 t
340.01 408.75 (1) 0.50 0.00 0.00 t
348.80 399.48 (1) 0.50 0.00 0.00 t
356.48 398.05 (1) 0.50 0.00 0.00 t
363.31 396.23 (1) 0.50 0.00 0.00 t
369.45 393.76 (1) 0.50 0.00 0.00 t
375.04 389.86 (1) 0.50 0.00 0.00 t
380.16 387.25 (1) 0.50 0.00 0.00 t
384.88 382.99 (1) 0.50 0.00 0.00 t
389.27 369.68 (1) 0.50 0.00 0.00 t
393.36 380.64 (1) 0.50 0.00 0.00 t
397.20 379.67 (1) 0.50 0.00 0.00 t
400.81 378.53 (1) 0.50 0.00 0.00 t
404.23 377.17 (1) 0.50 0.00 0.00 t
407.46 375.48 (1) 0.50 0.00 0.00 t
410.53 374.64 (1) 0.50 0.00 0.00 t
413.45 373.67 (1) 0.50 0.00 0.00 t
416.24 372.56 (1) 0.50 0.00 0.00 t
418.91 371.22 (1) 0.50 0.00 0.00 t
421.47 369.56 (1) 0.50 0.00 0.00 t
423.93 367.36 (1) 0.50 0.00 0.00 t
426.29 364.12 (1) 0.50 0.00 0.00 t
428.56 357.79 (1) 0.50 0.00 0.00 t
430.75 351.06 (1) 0.50 0.00 0.00 t
432.87 348.18 (1) 0.50 0.00 0.00 t
434.92 356.85 (1) 0.50 0.00 0.00 t
436.90 360.56 (1) 0.50 0.00 0.00 t
438.82 360.05 (1) 0.50 0.00 0.00 t
440.68 359.49 (1) 0.50 0.00 0.00 t
442.48 358.88 (1) 0.50 0.00 0.00 t
444.24 358.21 (1) 0.50 0.00 0.00 t
445.94 357.59 (1) 0.50 0.00 0.00 t
447.60 356.90 (1) 0.50 0.00 0.00 t
449.22 356.14 (1) 0.50 0.00 0.00 t
450.79 355.29 (1) 0.50 0.00 0.00 t
452.33 354.65 (1) 0.50 0.00 0.00 t
117.64 276.94 477.64 564.94 cl
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
np
192.53 344.26 m
432.69 344.26 l
o
np
192.53 344.26 m
192.53 337.66 l
o
np
248.78 344.26 m
248.78 337.66 l
o
np
291.33 344.26 m
291.33 337.66 l
o
np
333.88 344.26 m
333.88 337.66 l
o
np
390.13 344.26 m
390.13 337.66 l
o
np
432.69 344.26 m
432.69 337.66 l
o
/ps 11 def R 11 s
192.53 320.50 (20) 0.50 0.00 0.00 t
248.78 320.50 (50) 0.50 0.00 0.00 t
291.33 320.50 (100) 0.50 0.00 0.00 t
333.88 320.50 (200) 0.50 0.00 0.00 t
390.13 320.50 (500) 0.50 0.00 0.00 t
432.69 320.50 (1000) 0.50 0.00 0.00 t
np
171.76 349.67 m
171.76 539.93 l
o
np
171.76 349.67 m
165.16 349.67 l
o
np
171.76 397.24 m
165.16 397.24 l
o
np
171.76 444.80 m
165.16 444.80 l
o
np
171.76 492.37 m
165.16 492.37 l
o
np
171.76 539.93 m
165.16 539.93 l
o
155.92 349.67 (1e-11) 0.50 0.00 90.00 t
155.92 397.24 (1e-08) 0.50 0.00 90.00 t
155.92 444.80 (1e-05) 0.50 0.00 90.00 t
155.92 492.37 (1e-02) 0.50 0.00 90.00 t
155.92 539.93 (1e+01) 0.50 0.00 90.00 t
np
171.76 344.26 m
463.12 344.26 l
463.12 550.42 l
171.76 550.42 l
171.76 344.26 l
o
117.64 276.94 477.64 564.94 cl
/ps 11 def R 11 s
0.0000 0.0000 0.0000 rgb
317.44 294.10 (nombre d'�valuations) 0.50 0.00 0.00 t
129.52 447.34 (erreur) 0.50 0.00 90.00 t
171.76 344.26 463.12 550.42 cl
/ps 11 def R 11 s
1.0000 0.0000 0.0000 rgb
182.55 539.07 (2) 0.50 0.00 0.00 t
249.99 527.17 (2) 0.50 0.00 0.00 t
281.35 526.18 (2) 0.50 0.00 0.00 t
302.01 523.94 (2) 0.50 0.00 0.00 t
317.44 522.35 (2) 0.50 0.00 0.00 t
329.76 520.18 (2) 0.50 0.00 0.00 t
340.01 512.70 (2) 0.50 0.00 0.00 t
348.80 492.81 (2) 0.50 0.00 0.00 t
356.48 481.76 (2) 0.50 0.00 0.00 t
363.31 489.36 (2) 0.50 0.00 0.00 t
369.45 490.17 (2) 0.50 0.00 0.00 t
375.04 490.84 (2) 0.50 0.00 0.00 t
380.16 490.87 (2) 0.50 0.00 0.00 t
384.88 490.70 (2) 0.50 0.00 0.00 t
389.27 473.77 (2) 0.50 0.00 0.00 t
393.36 485.42 (2) 0.50 0.00 0.00 t
397.20 486.79 (2) 0.50 0.00 0.00 t
400.81 487.86 (2) 0.50 0.00 0.00 t
404.23 487.90 (2) 0.50 0.00 0.00 t
407.46 487.64 (2) 0.50 0.00 0.00 t
410.53 485.11 (2) 0.50 0.00 0.00 t
413.45 475.26 (2) 0.50 0.00 0.00 t
416.24 479.90 (2) 0.50 0.00 0.00 t
418.91 482.50 (2) 0.50 0.00 0.00 t
421.47 482.57 (2) 0.50 0.00 0.00 t
423.93 482.01 (2) 0.50 0.00 0.00 t
426.29 489.19 (2) 0.50 0.00 0.00 t
428.56 481.22 (2) 0.50 0.00 0.00 t
430.75 477.64 (2) 0.50 0.00 0.00 t
432.87 470.70 (2) 0.50 0.00 0.00 t
434.92 470.28 (2) 0.50 0.00 0.00 t
436.90 472.92 (2) 0.50 0.00 0.00 t
438.82 471.21 (2) 0.50 0.00 0.00 t
440.68 468.93 (2) 0.50 0.00 0.00 t
442.48 465.48 (2) 0.50 0.00 0.00 t
444.24 458.27 (2) 0.50 0.00 0.00 t
445.94 461.18 (2) 0.50 0.00 0.00 t
447.60 463.22 (2) 0.50 0.00 0.00 t
449.22 464.80 (2) 0.50 0.00 0.00 t
450.79 466.08 (2) 0.50 0.00 0.00 t
452.33 465.26 (2) 0.50 0.00 0.00 t
0.0000 0.0000 0.0000 rgb
0.75 setlinewidth
[] 0 setdash
349.99 543.98 443.32 504.38 r p1
359.89 527.06 (1) 0.50 0.00 0.00 t
1.0000 0.0000 0.0000 rgb
359.89 513.86 (2) 0.50 0.00 0.00 t
0.0000 0.0000 0.0000 rgb
374.74 527.08 (lisse) 0.00 0.00 0.00 t
374.74 513.90 (non-d�rivable) 0.00 0.00 0.00 t
ep
%%Trailer
%%Pages: 1
%%EOF
